module ibex_ex_block (alu_instr_first_cycle_i,
    branch_decision_o,
    clk_i,
    data_ind_timing_i,
    div_en_i,
    div_sel_i,
    ex_valid_o,
    mult_en_i,
    mult_sel_i,
    multdiv_ready_id_i,
    rst_ni,
    alu_adder_result_ex_o,
    alu_operand_a_i,
    alu_operand_b_i,
    alu_operator_i,
    branch_target_o,
    bt_a_operand_i,
    bt_b_operand_i,
    imd_val_d_o,
    imd_val_q_i,
    imd_val_we_o,
    multdiv_operand_a_i,
    multdiv_operand_b_i,
    multdiv_operator_i,
    multdiv_signed_mode_i,
    result_ex_o);
 input alu_instr_first_cycle_i;
 output branch_decision_o;
 input clk_i;
 input data_ind_timing_i;
 input div_en_i;
 input div_sel_i;
 output ex_valid_o;
 input mult_en_i;
 input mult_sel_i;
 input multdiv_ready_id_i;
 input rst_ni;
 output [31:0] alu_adder_result_ex_o;
 input [31:0] alu_operand_a_i;
 input [31:0] alu_operand_b_i;
 input [5:0] alu_operator_i;
 output [31:0] branch_target_o;
 input [31:0] bt_a_operand_i;
 input [31:0] bt_b_operand_i;
 output [67:0] imd_val_d_o;
 input [67:0] imd_val_q_i;
 output [1:0] imd_val_we_o;
 input [31:0] multdiv_operand_a_i;
 input [31:0] multdiv_operand_b_i;
 input [1:0] multdiv_operator_i;
 input [1:0] multdiv_signed_mode_i;
 output [31:0] result_ex_o;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire _3737_;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire _3747_;
 wire _3748_;
 wire _3749_;
 wire _3750_;
 wire _3751_;
 wire _3752_;
 wire _3753_;
 wire _3754_;
 wire _3755_;
 wire _3756_;
 wire _3757_;
 wire _3758_;
 wire _3759_;
 wire _3760_;
 wire _3761_;
 wire _3762_;
 wire _3763_;
 wire _3764_;
 wire _3765_;
 wire _3766_;
 wire _3767_;
 wire _3768_;
 wire _3769_;
 wire _3770_;
 wire _3771_;
 wire _3772_;
 wire _3773_;
 wire _3774_;
 wire _3775_;
 wire _3776_;
 wire _3777_;
 wire _3778_;
 wire _3779_;
 wire _3780_;
 wire _3781_;
 wire _3782_;
 wire _3783_;
 wire _3784_;
 wire _3785_;
 wire _3786_;
 wire _3787_;
 wire _3788_;
 wire _3789_;
 wire _3790_;
 wire _3791_;
 wire _3792_;
 wire _3793_;
 wire _3794_;
 wire _3795_;
 wire _3796_;
 wire _3797_;
 wire _3798_;
 wire _3799_;
 wire _3800_;
 wire _3801_;
 wire _3802_;
 wire _3803_;
 wire _3804_;
 wire _3805_;
 wire _3806_;
 wire _3807_;
 wire _3808_;
 wire _3809_;
 wire _3810_;
 wire _3811_;
 wire _3812_;
 wire _3813_;
 wire _3814_;
 wire _3815_;
 wire _3816_;
 wire _3817_;
 wire _3818_;
 wire _3819_;
 wire _3820_;
 wire _3821_;
 wire _3822_;
 wire _3823_;
 wire _3824_;
 wire _3825_;
 wire _3826_;
 wire _3827_;
 wire _3828_;
 wire _3829_;
 wire _3830_;
 wire _3831_;
 wire _3832_;
 wire _3833_;
 wire _3834_;
 wire _3835_;
 wire _3836_;
 wire _3837_;
 wire _3838_;
 wire _3839_;
 wire _3840_;
 wire _3841_;
 wire _3842_;
 wire _3843_;
 wire _3844_;
 wire _3845_;
 wire _3846_;
 wire _3847_;
 wire _3848_;
 wire _3849_;
 wire _3850_;
 wire _3851_;
 wire _3852_;
 wire _3853_;
 wire _3854_;
 wire _3855_;
 wire _3856_;
 wire _3857_;
 wire _3858_;
 wire _3859_;
 wire _3860_;
 wire _3861_;
 wire _3862_;
 wire _3863_;
 wire _3864_;
 wire _3865_;
 wire _3866_;
 wire _3867_;
 wire _3868_;
 wire _3869_;
 wire _3870_;
 wire _3871_;
 wire _3872_;
 wire _3873_;
 wire _3874_;
 wire _3875_;
 wire _3876_;
 wire _3877_;
 wire _3878_;
 wire _3879_;
 wire _3880_;
 wire _3881_;
 wire _3882_;
 wire _3883_;
 wire _3884_;
 wire _3885_;
 wire _3886_;
 wire _3887_;
 wire _3888_;
 wire _3889_;
 wire _3890_;
 wire _3891_;
 wire _3892_;
 wire _3893_;
 wire _3894_;
 wire _3895_;
 wire _3896_;
 wire _3897_;
 wire _3898_;
 wire _3899_;
 wire _3900_;
 wire _3901_;
 wire _3902_;
 wire _3903_;
 wire _3904_;
 wire _3905_;
 wire _3906_;
 wire _3907_;
 wire _3908_;
 wire _3909_;
 wire _3910_;
 wire _3911_;
 wire _3912_;
 wire _3913_;
 wire _3914_;
 wire _3915_;
 wire _3916_;
 wire _3917_;
 wire _3918_;
 wire _3919_;
 wire _3920_;
 wire _3921_;
 wire _3922_;
 wire _3923_;
 wire _3924_;
 wire _3925_;
 wire _3926_;
 wire _3927_;
 wire _3928_;
 wire _3929_;
 wire _3930_;
 wire _3931_;
 wire _3932_;
 wire _3933_;
 wire _3934_;
 wire _3935_;
 wire _3936_;
 wire _3937_;
 wire _3938_;
 wire _3939_;
 wire _3940_;
 wire _3941_;
 wire _3942_;
 wire _3943_;
 wire _3944_;
 wire _3945_;
 wire _3946_;
 wire _3947_;
 wire _3948_;
 wire _3949_;
 wire _3950_;
 wire _3951_;
 wire _3952_;
 wire _3953_;
 wire _3954_;
 wire _3955_;
 wire _3956_;
 wire _3957_;
 wire _3958_;
 wire _3959_;
 wire _3960_;
 wire _3961_;
 wire _3962_;
 wire _3963_;
 wire _3964_;
 wire _3965_;
 wire _3966_;
 wire _3967_;
 wire _3968_;
 wire _3969_;
 wire _3970_;
 wire _3971_;
 wire _3972_;
 wire _3973_;
 wire _3974_;
 wire _3975_;
 wire _3976_;
 wire _3977_;
 wire _3978_;
 wire _3979_;
 wire _3980_;
 wire _3981_;
 wire _3982_;
 wire _3983_;
 wire _3984_;
 wire _3985_;
 wire _3986_;
 wire _3987_;
 wire _3988_;
 wire _3989_;
 wire _3990_;
 wire _3991_;
 wire _3992_;
 wire _3993_;
 wire _3994_;
 wire _3995_;
 wire _3996_;
 wire _3997_;
 wire _3998_;
 wire _3999_;
 wire _4000_;
 wire _4001_;
 wire _4002_;
 wire _4003_;
 wire _4004_;
 wire _4005_;
 wire _4006_;
 wire _4007_;
 wire _4008_;
 wire _4009_;
 wire _4010_;
 wire _4011_;
 wire _4012_;
 wire _4013_;
 wire _4014_;
 wire _4015_;
 wire _4016_;
 wire _4017_;
 wire _4018_;
 wire _4019_;
 wire _4020_;
 wire _4021_;
 wire _4022_;
 wire _4023_;
 wire _4024_;
 wire _4025_;
 wire _4026_;
 wire _4027_;
 wire _4028_;
 wire _4029_;
 wire _4030_;
 wire _4031_;
 wire _4032_;
 wire _4033_;
 wire _4034_;
 wire _4035_;
 wire _4036_;
 wire _4037_;
 wire _4038_;
 wire _4039_;
 wire _4040_;
 wire _4041_;
 wire _4042_;
 wire _4043_;
 wire _4044_;
 wire _4045_;
 wire _4046_;
 wire _4047_;
 wire _4048_;
 wire _4049_;
 wire _4050_;
 wire _4051_;
 wire _4052_;
 wire _4053_;
 wire _4054_;
 wire _4055_;
 wire _4056_;
 wire _4057_;
 wire _4058_;
 wire _4059_;
 wire _4060_;
 wire _4061_;
 wire _4062_;
 wire _4063_;
 wire _4064_;
 wire _4065_;
 wire _4066_;
 wire _4067_;
 wire _4068_;
 wire _4069_;
 wire _4070_;
 wire _4071_;
 wire _4072_;
 wire _4073_;
 wire _4074_;
 wire _4075_;
 wire _4076_;
 wire _4077_;
 wire _4078_;
 wire _4079_;
 wire _4080_;
 wire _4081_;
 wire _4082_;
 wire _4083_;
 wire _4084_;
 wire _4085_;
 wire _4086_;
 wire _4087_;
 wire _4088_;
 wire _4089_;
 wire _4090_;
 wire _4091_;
 wire _4092_;
 wire _4093_;
 wire _4094_;
 wire _4095_;
 wire _4096_;
 wire _4097_;
 wire _4098_;
 wire _4099_;
 wire _4100_;
 wire _4101_;
 wire _4102_;
 wire _4103_;
 wire _4104_;
 wire _4105_;
 wire _4106_;
 wire _4107_;
 wire _4108_;
 wire _4109_;
 wire _4110_;
 wire _4111_;
 wire _4112_;
 wire _4113_;
 wire _4114_;
 wire _4115_;
 wire _4116_;
 wire _4117_;
 wire _4118_;
 wire _4119_;
 wire _4120_;
 wire clknet_0_clk_i;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire \genblk3.gen_multdiv_fast.multdiv_i.div_by_zero_q ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[2] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[3] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[4] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.div_valid ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[1] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[2] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.md_state_q[0] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.md_state_q[2] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.md_state_q[5] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.md_state_q[6] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[0] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[10] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[11] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[12] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[13] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[14] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[15] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[16] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[17] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[18] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[19] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[1] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[20] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[21] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[22] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[23] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[24] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[25] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[26] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[27] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[28] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[29] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[2] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[30] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[31] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[3] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[4] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[5] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[6] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[7] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[8] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[9] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[0] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[10] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[11] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[12] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[13] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[14] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[15] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[16] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[17] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[18] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[19] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[1] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[20] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[21] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[22] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[23] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[24] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[25] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[26] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[27] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[28] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[29] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[2] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[30] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[31] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[3] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[4] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[5] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[6] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[7] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[8] ;
 wire \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[9] ;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire clknet_3_0_0_clk_i;
 wire clknet_3_1_0_clk_i;
 wire clknet_3_2_0_clk_i;
 wire clknet_3_3_0_clk_i;
 wire clknet_3_4_0_clk_i;
 wire clknet_3_5_0_clk_i;
 wire clknet_3_6_0_clk_i;
 wire clknet_3_7_0_clk_i;
 wire net365;
 wire net366;

 sky130_fd_sc_hs__clkbuf_8 _4122_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3] ),
    .X(_0081_));
 sky130_fd_sc_hs__nand2_1 _4123_ (.A(net187),
    .B(net120),
    .Y(_0082_));
 sky130_fd_sc_hs__nor2_8 _4124_ (.A(net185),
    .B(net186),
    .Y(_0083_));
 sky130_fd_sc_hs__clkbuf_8 _4125_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[1] ),
    .X(_0084_));
 sky130_fd_sc_hs__nor2b_4 _4126_ (.A(_0083_),
    .B_N(_0084_),
    .Y(_0085_));
 sky130_fd_sc_hs__clkbuf_8 _4127_ (.A(_0085_),
    .X(_0086_));
 sky130_fd_sc_hs__a21oi_4 _4128_ (.A1(_0084_),
    .A2(_0083_),
    .B1(_0081_),
    .Y(_0087_));
 sky130_fd_sc_hs__o21ai_4 _4129_ (.A1(net187),
    .A2(_0087_),
    .B1(net120),
    .Y(_0088_));
 sky130_fd_sc_hs__inv_1 _4130_ (.A(_0088_),
    .Y(_0089_));
 sky130_fd_sc_hs__a22o_1 _4131_ (.A1(_0081_),
    .A2(_0082_),
    .B1(_0086_),
    .B2(_0089_),
    .X(_0001_));
 sky130_fd_sc_hs__buf_8 _4132_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.md_state_q[2] ),
    .X(_0090_));
 sky130_fd_sc_hs__clkbuf_16 _4133_ (.A(_0090_),
    .X(_0091_));
 sky130_fd_sc_hs__inv_2 _4134_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.div_valid ),
    .Y(_0092_));
 sky130_fd_sc_hs__o21a_1 _4135_ (.A1(_0092_),
    .A2(net187),
    .B1(net79),
    .X(_0093_));
 sky130_fd_sc_hs__clkbuf_8 _4136_ (.A(_0093_),
    .X(_0094_));
 sky130_fd_sc_hs__buf_8 _4137_ (.A(_3710_),
    .X(_0095_));
 sky130_fd_sc_hs__clkbuf_8 _4138_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[4] ),
    .X(_0096_));
 sky130_fd_sc_hs__buf_8 _4139_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .X(_0097_));
 sky130_fd_sc_hs__clkbuf_8 _4140_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .X(_0098_));
 sky130_fd_sc_hs__nor3_4 _4141_ (.A(_0096_),
    .B(_0097_),
    .C(_0098_),
    .Y(_0099_));
 sky130_fd_sc_hs__and2_1 _4142_ (.A(_0095_),
    .B(_0099_),
    .X(_0100_));
 sky130_fd_sc_hs__nand2_1 _4143_ (.A(_0094_),
    .B(_0100_),
    .Y(_0101_));
 sky130_fd_sc_hs__buf_8 _4144_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .X(_0102_));
 sky130_fd_sc_hs__buf_8 _4145_ (.A(_0102_),
    .X(_0103_));
 sky130_fd_sc_hs__a22o_1 _4146_ (.A1(_0091_),
    .A2(_0094_),
    .B1(_0101_),
    .B2(_0103_),
    .X(_0005_));
 sky130_fd_sc_hs__inv_1 _4147_ (.A(net2),
    .Y(_3937_));
 sky130_fd_sc_hs__inv_1 _4148_ (.A(net21),
    .Y(_3942_));
 sky130_fd_sc_hs__inv_1 _4149_ (.A(net32),
    .Y(_3947_));
 sky130_fd_sc_hs__buf_8 _4150_ (.A(mult_sel_i),
    .X(_0104_));
 sky130_fd_sc_hs__buf_8 _4151_ (.A(net80),
    .X(_0105_));
 sky130_fd_sc_hs__nor2_4 _4152_ (.A(_0104_),
    .B(_0105_),
    .Y(_0106_));
 sky130_fd_sc_hs__buf_8 _4153_ (.A(_0106_),
    .X(_0107_));
 sky130_fd_sc_hs__buf_4 _4154_ (.A(_0107_),
    .X(_0108_));
 sky130_fd_sc_hs__buf_16 _4155_ (.A(_0108_),
    .X(_0109_));
 sky130_fd_sc_hs__clkbuf_8 _4156_ (.A(alu_operator_i[2]),
    .X(_0110_));
 sky130_fd_sc_hs__and3_4 _4157_ (.A(_0110_),
    .B(net77),
    .C(_3569_),
    .X(_0111_));
 sky130_fd_sc_hs__buf_4 _4158_ (.A(_3572_),
    .X(_0112_));
 sky130_fd_sc_hs__nor3b_4 _4159_ (.A(_0110_),
    .B(net77),
    .C_N(_0112_),
    .Y(_0113_));
 sky130_fd_sc_hs__buf_4 _4160_ (.A(alu_operator_i[3]),
    .X(_0114_));
 sky130_fd_sc_hs__nor2_4 _4161_ (.A(_0114_),
    .B(net76),
    .Y(_0115_));
 sky130_fd_sc_hs__o21ai_4 _4162_ (.A1(_0111_),
    .A2(_0113_),
    .B1(_0115_),
    .Y(_0116_));
 sky130_fd_sc_hs__nor2b_4 _4163_ (.A(net77),
    .B_N(net76),
    .Y(_0117_));
 sky130_fd_sc_hs__buf_4 _4164_ (.A(_3568_),
    .X(_0118_));
 sky130_fd_sc_hs__nand3b_2 _4165_ (.A_N(_0118_),
    .B(_0114_),
    .C(_0110_),
    .Y(_0119_));
 sky130_fd_sc_hs__or3_2 _4166_ (.A(_0110_),
    .B(_0114_),
    .C(_3574_),
    .X(_0120_));
 sky130_fd_sc_hs__nand3_4 _4167_ (.A(_0117_),
    .B(_0119_),
    .C(_0120_),
    .Y(_0121_));
 sky130_fd_sc_hs__nand3_2 _4168_ (.A(_0109_),
    .B(_0116_),
    .C(_0121_),
    .Y(_2226_));
 sky130_fd_sc_hs__inv_1 _4169_ (.A(net35),
    .Y(_3953_));
 sky130_fd_sc_hs__inv_1 _4170_ (.A(net36),
    .Y(_3959_));
 sky130_fd_sc_hs__inv_1 _4171_ (.A(net37),
    .Y(_3965_));
 sky130_fd_sc_hs__inv_1 _4172_ (.A(net38),
    .Y(_3971_));
 sky130_fd_sc_hs__inv_1 _4173_ (.A(net39),
    .Y(_3977_));
 sky130_fd_sc_hs__inv_1 _4174_ (.A(net40),
    .Y(_3983_));
 sky130_fd_sc_hs__inv_1 _4175_ (.A(net41),
    .Y(_3989_));
 sky130_fd_sc_hs__inv_1 _4176_ (.A(net3),
    .Y(_3995_));
 sky130_fd_sc_hs__inv_1 _4177_ (.A(net4),
    .Y(_4001_));
 sky130_fd_sc_hs__inv_1 _4178_ (.A(net5),
    .Y(_4007_));
 sky130_fd_sc_hs__inv_1 _4179_ (.A(net6),
    .Y(_4013_));
 sky130_fd_sc_hs__inv_1 _4180_ (.A(net7),
    .Y(_4019_));
 sky130_fd_sc_hs__inv_2 _4181_ (.A(net8),
    .Y(_4025_));
 sky130_fd_sc_hs__clkinv_2 _4182_ (.A(net17),
    .Y(_4031_));
 sky130_fd_sc_hs__inv_1 _4183_ (.A(net18),
    .Y(_4037_));
 sky130_fd_sc_hs__inv_1 _4184_ (.A(net19),
    .Y(_4043_));
 sky130_fd_sc_hs__inv_1 _4185_ (.A(net20),
    .Y(_4049_));
 sky130_fd_sc_hs__inv_1 _4186_ (.A(net22),
    .Y(_4055_));
 sky130_fd_sc_hs__inv_1 _4187_ (.A(net23),
    .Y(_4061_));
 sky130_fd_sc_hs__inv_1 _4188_ (.A(net24),
    .Y(_4067_));
 sky130_fd_sc_hs__inv_1 _4189_ (.A(net25),
    .Y(_4073_));
 sky130_fd_sc_hs__inv_1 _4190_ (.A(net26),
    .Y(_4079_));
 sky130_fd_sc_hs__inv_1 _4191_ (.A(net27),
    .Y(_4085_));
 sky130_fd_sc_hs__inv_1 _4192_ (.A(net28),
    .Y(_4091_));
 sky130_fd_sc_hs__inv_1 _4193_ (.A(net29),
    .Y(_4097_));
 sky130_fd_sc_hs__inv_1 _4194_ (.A(net30),
    .Y(_4103_));
 sky130_fd_sc_hs__inv_1 _4195_ (.A(net31),
    .Y(_4109_));
 sky130_fd_sc_hs__inv_1 _4196_ (.A(net33),
    .Y(_4115_));
 sky130_fd_sc_hs__inv_2 _4197_ (.A(net34),
    .Y(_3927_));
 sky130_fd_sc_hs__clkbuf_16 _4198_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.md_state_q[0] ),
    .X(_0122_));
 sky130_fd_sc_hs__buf_8 _4199_ (.A(_0122_),
    .X(_0123_));
 sky130_fd_sc_hs__and2_2 _4200_ (.A(_3657_),
    .B(_3661_),
    .X(_0124_));
 sky130_fd_sc_hs__nand2_4 _4201_ (.A(_3669_),
    .B(_3673_),
    .Y(_0125_));
 sky130_fd_sc_hs__buf_4 _4202_ (.A(_3665_),
    .X(_0126_));
 sky130_fd_sc_hs__nand2_2 _4203_ (.A(_0126_),
    .B(_3677_),
    .Y(_0127_));
 sky130_fd_sc_hs__clkbuf_8 _4204_ (.A(_3681_),
    .X(_0128_));
 sky130_fd_sc_hs__nand2_2 _4205_ (.A(_0128_),
    .B(_3685_),
    .Y(_0129_));
 sky130_fd_sc_hs__nor3_4 _4206_ (.A(_0125_),
    .B(_0127_),
    .C(_0129_),
    .Y(_0130_));
 sky130_fd_sc_hs__nand2_1 _4207_ (.A(_0124_),
    .B(_0130_),
    .Y(_0131_));
 sky130_fd_sc_hs__or2_4 _4208_ (.A(_0104_),
    .B(net80),
    .X(_0132_));
 sky130_fd_sc_hs__o21a_2 _4209_ (.A1(_0111_),
    .A2(_0113_),
    .B1(_0115_),
    .X(_0133_));
 sky130_fd_sc_hs__and3_2 _4210_ (.A(_0117_),
    .B(_0119_),
    .C(_0120_),
    .X(_0134_));
 sky130_fd_sc_hs__and2_2 _4211_ (.A(_3581_),
    .B(_3577_),
    .X(_0135_));
 sky130_fd_sc_hs__o31ai_4 _4212_ (.A1(_0132_),
    .A2(_0133_),
    .A3(_0134_),
    .B1(_0135_),
    .Y(_0136_));
 sky130_fd_sc_hs__inv_4 _4213_ (.A(_3588_),
    .Y(_0137_));
 sky130_fd_sc_hs__o21ai_4 _4214_ (.A1(_3585_),
    .A2(_3584_),
    .B1(_3589_),
    .Y(_0138_));
 sky130_fd_sc_hs__nand2_8 _4215_ (.A(_3593_),
    .B(_3597_),
    .Y(_0139_));
 sky130_fd_sc_hs__a21oi_4 _4216_ (.A1(_0137_),
    .A2(_0138_),
    .B1(_0139_),
    .Y(_0140_));
 sky130_fd_sc_hs__nand2_4 _4217_ (.A(_3601_),
    .B(_0140_),
    .Y(_0141_));
 sky130_fd_sc_hs__a21o_4 _4218_ (.A1(_3597_),
    .A2(_3592_),
    .B1(_3596_),
    .X(_0142_));
 sky130_fd_sc_hs__a21oi_4 _4219_ (.A1(_3581_),
    .A2(_3576_),
    .B1(_3580_),
    .Y(_0143_));
 sky130_fd_sc_hs__a21oi_2 _4220_ (.A1(_3589_),
    .A2(_3584_),
    .B1(_3588_),
    .Y(_0144_));
 sky130_fd_sc_hs__a221oi_2 _4221_ (.A1(_0137_),
    .A2(_0138_),
    .B1(_0143_),
    .B2(_0144_),
    .C1(_0139_),
    .Y(_0145_));
 sky130_fd_sc_hs__o21ai_2 _4222_ (.A1(_0142_),
    .A2(_0145_),
    .B1(_3601_),
    .Y(_0146_));
 sky130_fd_sc_hs__o21ai_4 _4223_ (.A1(_0136_),
    .A2(_0141_),
    .B1(_0146_),
    .Y(_0147_));
 sky130_fd_sc_hs__and2_1 _4224_ (.A(_3605_),
    .B(_3609_),
    .X(_0148_));
 sky130_fd_sc_hs__clkbuf_8 _4225_ (.A(_3633_),
    .X(_0149_));
 sky130_fd_sc_hs__inv_2 _4226_ (.A(_3625_),
    .Y(_0150_));
 sky130_fd_sc_hs__inv_2 _4227_ (.A(_3629_),
    .Y(_0151_));
 sky130_fd_sc_hs__nor2_8 _4228_ (.A(_0150_),
    .B(_0151_),
    .Y(_0152_));
 sky130_fd_sc_hs__nand2_8 _4229_ (.A(_0149_),
    .B(_0152_),
    .Y(_0153_));
 sky130_fd_sc_hs__clkbuf_8 _4230_ (.A(_3617_),
    .X(_0154_));
 sky130_fd_sc_hs__nand3_4 _4231_ (.A(_3613_),
    .B(_0154_),
    .C(_3621_),
    .Y(_0155_));
 sky130_fd_sc_hs__nor2_4 _4232_ (.A(_0153_),
    .B(_0155_),
    .Y(_0156_));
 sky130_fd_sc_hs__inv_2 _4233_ (.A(_3609_),
    .Y(_0157_));
 sky130_fd_sc_hs__a21oi_1 _4234_ (.A1(_3605_),
    .A2(_3600_),
    .B1(_3604_),
    .Y(_0158_));
 sky130_fd_sc_hs__o21ba_4 _4235_ (.A1(_0157_),
    .A2(_0158_),
    .B1_N(_3608_),
    .X(_0159_));
 sky130_fd_sc_hs__a21o_1 _4236_ (.A1(_0154_),
    .A2(_3612_),
    .B1(_3616_),
    .X(_0160_));
 sky130_fd_sc_hs__a21oi_4 _4237_ (.A1(_3621_),
    .A2(_0160_),
    .B1(_3620_),
    .Y(_0161_));
 sky130_fd_sc_hs__o21ai_4 _4238_ (.A1(_0159_),
    .A2(_0155_),
    .B1(_0161_),
    .Y(_0162_));
 sky130_fd_sc_hs__and3_4 _4239_ (.A(_3625_),
    .B(_3629_),
    .C(_0149_),
    .X(_0163_));
 sky130_fd_sc_hs__a32oi_4 _4240_ (.A1(_0147_),
    .A2(_0148_),
    .A3(_0156_),
    .B1(_0162_),
    .B2(_0163_),
    .Y(_0164_));
 sky130_fd_sc_hs__a21o_2 _4241_ (.A1(_3629_),
    .A2(_3624_),
    .B1(_3628_),
    .X(_0165_));
 sky130_fd_sc_hs__a21o_2 _4242_ (.A1(_0149_),
    .A2(_0165_),
    .B1(_3632_),
    .X(_0166_));
 sky130_fd_sc_hs__buf_4 _4243_ (.A(_3653_),
    .X(_0167_));
 sky130_fd_sc_hs__clkbuf_8 _4244_ (.A(_3649_),
    .X(_0168_));
 sky130_fd_sc_hs__inv_2 _4245_ (.A(_0168_),
    .Y(_0169_));
 sky130_fd_sc_hs__a21oi_2 _4246_ (.A1(_3645_),
    .A2(_3640_),
    .B1(_3644_),
    .Y(_0170_));
 sky130_fd_sc_hs__o21bai_1 _4247_ (.A1(_0169_),
    .A2(_0170_),
    .B1_N(_3648_),
    .Y(_0171_));
 sky130_fd_sc_hs__a21oi_1 _4248_ (.A1(_0167_),
    .A2(_0171_),
    .B1(_3652_),
    .Y(_0172_));
 sky130_fd_sc_hs__nor3b_4 _4249_ (.A(_3636_),
    .B(_0166_),
    .C_N(_0172_),
    .Y(_0173_));
 sky130_fd_sc_hs__inv_1 _4250_ (.A(_0167_),
    .Y(_0174_));
 sky130_fd_sc_hs__clkbuf_4 _4251_ (.A(_3641_),
    .X(_0175_));
 sky130_fd_sc_hs__nand2_1 _4252_ (.A(_0175_),
    .B(_3645_),
    .Y(_0176_));
 sky130_fd_sc_hs__clkbuf_4 _4253_ (.A(_3637_),
    .X(_0177_));
 sky130_fd_sc_hs__nor2_1 _4254_ (.A(_0177_),
    .B(_3636_),
    .Y(_0178_));
 sky130_fd_sc_hs__o41a_2 _4255_ (.A1(_0169_),
    .A2(_0174_),
    .A3(_0176_),
    .A4(_0178_),
    .B1(_0172_),
    .X(_0179_));
 sky130_fd_sc_hs__a21o_4 _4256_ (.A1(_0164_),
    .A2(_0173_),
    .B1(_0179_),
    .X(_0180_));
 sky130_fd_sc_hs__inv_2 _4257_ (.A(_3673_),
    .Y(_0181_));
 sky130_fd_sc_hs__inv_1 _4258_ (.A(_3677_),
    .Y(_0182_));
 sky130_fd_sc_hs__a21o_1 _4259_ (.A1(_3661_),
    .A2(_3656_),
    .B1(_3660_),
    .X(_0183_));
 sky130_fd_sc_hs__a21o_1 _4260_ (.A1(_0126_),
    .A2(_0183_),
    .B1(_3664_),
    .X(_0184_));
 sky130_fd_sc_hs__a21oi_4 _4261_ (.A1(_3669_),
    .A2(_0184_),
    .B1(_3668_),
    .Y(_0185_));
 sky130_fd_sc_hs__a21oi_1 _4262_ (.A1(_3677_),
    .A2(_3672_),
    .B1(_3676_),
    .Y(_0186_));
 sky130_fd_sc_hs__o31a_1 _4263_ (.A1(_0181_),
    .A2(_0182_),
    .A3(_0185_),
    .B1(_0186_),
    .X(_0187_));
 sky130_fd_sc_hs__a21oi_2 _4264_ (.A1(_3685_),
    .A2(_3680_),
    .B1(_3684_),
    .Y(_0188_));
 sky130_fd_sc_hs__o21a_1 _4265_ (.A1(_0129_),
    .A2(_0187_),
    .B1(_0188_),
    .X(_0189_));
 sky130_fd_sc_hs__nor2_1 _4266_ (.A(_3688_),
    .B(_3692_),
    .Y(_0190_));
 sky130_fd_sc_hs__o211a_1 _4267_ (.A1(_0131_),
    .A2(_0180_),
    .B1(_0189_),
    .C1(_0190_),
    .X(_0191_));
 sky130_fd_sc_hs__buf_2 _4268_ (.A(_3689_),
    .X(_0192_));
 sky130_fd_sc_hs__or2_1 _4269_ (.A(_0192_),
    .B(_3688_),
    .X(_0193_));
 sky130_fd_sc_hs__a21oi_2 _4270_ (.A1(_3693_),
    .A2(_0193_),
    .B1(_3692_),
    .Y(_0194_));
 sky130_fd_sc_hs__nor3_4 _4271_ (.A(_3697_),
    .B(_0191_),
    .C(_0194_),
    .Y(_0195_));
 sky130_fd_sc_hs__o21a_2 _4272_ (.A1(_0191_),
    .A2(_0194_),
    .B1(_3697_),
    .X(_0196_));
 sky130_fd_sc_hs__or2_1 _4273_ (.A(_0195_),
    .B(_0196_),
    .X(_0197_));
 sky130_fd_sc_hs__clkbuf_16 _4274_ (.A(_0197_),
    .X(net214));
 sky130_fd_sc_hs__a21oi_1 _4275_ (.A1(_3669_),
    .A2(_3664_),
    .B1(_3668_),
    .Y(_0198_));
 sky130_fd_sc_hs__o21bai_1 _4276_ (.A1(_0181_),
    .A2(_0198_),
    .B1_N(_3672_),
    .Y(_0199_));
 sky130_fd_sc_hs__nand2_8 _4277_ (.A(_3605_),
    .B(_3609_),
    .Y(_0200_));
 sky130_fd_sc_hs__nor2_2 _4278_ (.A(_0155_),
    .B(_0200_),
    .Y(_0201_));
 sky130_fd_sc_hs__a21o_1 _4279_ (.A1(_0152_),
    .A2(_0162_),
    .B1(_0165_),
    .X(_0202_));
 sky130_fd_sc_hs__a31oi_4 _4280_ (.A1(_0152_),
    .A2(_0147_),
    .A3(_0201_),
    .B1(_0202_),
    .Y(_0203_));
 sky130_fd_sc_hs__nand4_2 _4281_ (.A(_0149_),
    .B(_0177_),
    .C(_0175_),
    .D(_3645_),
    .Y(_0204_));
 sky130_fd_sc_hs__nand3_2 _4282_ (.A(_0168_),
    .B(_0167_),
    .C(_0124_),
    .Y(_0205_));
 sky130_fd_sc_hs__a21oi_2 _4283_ (.A1(_0177_),
    .A2(_3632_),
    .B1(_3636_),
    .Y(_0206_));
 sky130_fd_sc_hs__o21ai_4 _4284_ (.A1(_0176_),
    .A2(_0206_),
    .B1(_0170_),
    .Y(_0207_));
 sky130_fd_sc_hs__a21oi_1 _4285_ (.A1(_0168_),
    .A2(_0207_),
    .B1(_3648_),
    .Y(_0208_));
 sky130_fd_sc_hs__o21bai_1 _4286_ (.A1(_0174_),
    .A2(_0208_),
    .B1_N(_3652_),
    .Y(_0209_));
 sky130_fd_sc_hs__a21oi_2 _4287_ (.A1(_0124_),
    .A2(_0209_),
    .B1(_0183_),
    .Y(_0210_));
 sky130_fd_sc_hs__o31ai_4 _4288_ (.A1(_0203_),
    .A2(_0204_),
    .A3(_0205_),
    .B1(_0210_),
    .Y(_0211_));
 sky130_fd_sc_hs__nor2_2 _4289_ (.A(_0125_),
    .B(_0127_),
    .Y(_0212_));
 sky130_fd_sc_hs__a221oi_4 _4290_ (.A1(_3677_),
    .A2(_0199_),
    .B1(_0211_),
    .B2(_0212_),
    .C1(_3676_),
    .Y(_0213_));
 sky130_fd_sc_hs__xnor2_4 _4291_ (.A(_0128_),
    .B(_0213_),
    .Y(net209));
 sky130_fd_sc_hs__a21o_1 _4292_ (.A1(_3673_),
    .A2(_3668_),
    .B1(_3672_),
    .X(_0214_));
 sky130_fd_sc_hs__a21oi_2 _4293_ (.A1(_3657_),
    .A2(_3652_),
    .B1(_3656_),
    .Y(_0215_));
 sky130_fd_sc_hs__nand2_1 _4294_ (.A(_3661_),
    .B(_0126_),
    .Y(_0216_));
 sky130_fd_sc_hs__a21oi_1 _4295_ (.A1(_0126_),
    .A2(_3660_),
    .B1(_3664_),
    .Y(_0217_));
 sky130_fd_sc_hs__o21ai_4 _4296_ (.A1(_0215_),
    .A2(_0216_),
    .B1(_0217_),
    .Y(_0218_));
 sky130_fd_sc_hs__and4_2 _4297_ (.A(_0167_),
    .B(_3657_),
    .C(_3661_),
    .D(_0126_),
    .X(_0219_));
 sky130_fd_sc_hs__a21oi_4 _4298_ (.A1(_0175_),
    .A2(_3636_),
    .B1(_3640_),
    .Y(_0220_));
 sky130_fd_sc_hs__nand2_2 _4299_ (.A(_3645_),
    .B(_0168_),
    .Y(_0221_));
 sky130_fd_sc_hs__a21oi_4 _4300_ (.A1(_0168_),
    .A2(_3644_),
    .B1(_3648_),
    .Y(_0222_));
 sky130_fd_sc_hs__o21ai_4 _4301_ (.A1(_0220_),
    .A2(_0221_),
    .B1(_0222_),
    .Y(_0223_));
 sky130_fd_sc_hs__a21oi_1 _4302_ (.A1(_3625_),
    .A2(_3620_),
    .B1(_3624_),
    .Y(_0224_));
 sky130_fd_sc_hs__nand2_1 _4303_ (.A(_3629_),
    .B(_0149_),
    .Y(_0225_));
 sky130_fd_sc_hs__a21oi_1 _4304_ (.A1(_0149_),
    .A2(_3628_),
    .B1(_3632_),
    .Y(_0226_));
 sky130_fd_sc_hs__o21ai_2 _4305_ (.A1(_0224_),
    .A2(_0225_),
    .B1(_0226_),
    .Y(_0227_));
 sky130_fd_sc_hs__and4_1 _4306_ (.A(_0177_),
    .B(_0175_),
    .C(_3645_),
    .D(_0168_),
    .X(_0228_));
 sky130_fd_sc_hs__and2_1 _4307_ (.A(_0219_),
    .B(_0228_),
    .X(_0229_));
 sky130_fd_sc_hs__a22oi_4 _4308_ (.A1(_0219_),
    .A2(_0223_),
    .B1(_0227_),
    .B2(_0229_),
    .Y(_0230_));
 sky130_fd_sc_hs__nor2b_4 _4309_ (.A(_0218_),
    .B_N(_0230_),
    .Y(_0231_));
 sky130_fd_sc_hs__nand2_1 _4310_ (.A(_3613_),
    .B(_0154_),
    .Y(_0232_));
 sky130_fd_sc_hs__inv_2 _4311_ (.A(_0232_),
    .Y(_0233_));
 sky130_fd_sc_hs__and4_2 _4312_ (.A(_3621_),
    .B(_0163_),
    .C(_0219_),
    .D(_0228_),
    .X(_0234_));
 sky130_fd_sc_hs__a211oi_4 _4313_ (.A1(_3581_),
    .A2(_2229_),
    .B1(_3580_),
    .C1(_3584_),
    .Y(_0235_));
 sky130_fd_sc_hs__nor3_4 _4314_ (.A(_0138_),
    .B(_0139_),
    .C(_0235_),
    .Y(_0236_));
 sky130_fd_sc_hs__o21bai_4 _4315_ (.A1(_0137_),
    .A2(_0139_),
    .B1_N(_0142_),
    .Y(_0237_));
 sky130_fd_sc_hs__a21oi_4 _4316_ (.A1(_3609_),
    .A2(_3604_),
    .B1(_3608_),
    .Y(_0238_));
 sky130_fd_sc_hs__or4b_1 _4317_ (.A(_3600_),
    .B(_0236_),
    .C(_0237_),
    .D_N(_0238_),
    .X(_0239_));
 sky130_fd_sc_hs__clkbuf_4 _4318_ (.A(_0239_),
    .X(_0240_));
 sky130_fd_sc_hs__nor2_2 _4319_ (.A(_3601_),
    .B(_3600_),
    .Y(_0241_));
 sky130_fd_sc_hs__o21ai_4 _4320_ (.A1(_0200_),
    .A2(_0241_),
    .B1(_0238_),
    .Y(_0242_));
 sky130_fd_sc_hs__nand4_2 _4321_ (.A(_0233_),
    .B(_0234_),
    .C(_0240_),
    .D(_0242_),
    .Y(_0243_));
 sky130_fd_sc_hs__and2_1 _4322_ (.A(_0154_),
    .B(_3612_),
    .X(_0244_));
 sky130_fd_sc_hs__o21ai_4 _4323_ (.A1(_3616_),
    .A2(_0244_),
    .B1(_0234_),
    .Y(_0245_));
 sky130_fd_sc_hs__a31oi_4 _4324_ (.A1(_0231_),
    .A2(_0243_),
    .A3(_0245_),
    .B1(_0125_),
    .Y(_0246_));
 sky130_fd_sc_hs__o21ai_4 _4325_ (.A1(_0214_),
    .A2(_0246_),
    .B1(_3677_),
    .Y(_0247_));
 sky130_fd_sc_hs__or3_2 _4326_ (.A(_3677_),
    .B(_0214_),
    .C(_0246_),
    .X(_0248_));
 sky130_fd_sc_hs__and2_4 _4327_ (.A(_0247_),
    .B(_0248_),
    .X(net208));
 sky130_fd_sc_hs__nand4_2 _4328_ (.A(_0126_),
    .B(_3669_),
    .C(_3673_),
    .D(_0124_),
    .Y(_0249_));
 sky130_fd_sc_hs__a211oi_4 _4329_ (.A1(_0164_),
    .A2(_0173_),
    .B1(_0179_),
    .C1(_0249_),
    .Y(_0250_));
 sky130_fd_sc_hs__a21oi_1 _4330_ (.A1(_0126_),
    .A2(_3669_),
    .B1(_3673_),
    .Y(_0251_));
 sky130_fd_sc_hs__nand2_1 _4331_ (.A(_0185_),
    .B(_0251_),
    .Y(_0252_));
 sky130_fd_sc_hs__nor2_1 _4332_ (.A(_3673_),
    .B(_0124_),
    .Y(_0253_));
 sky130_fd_sc_hs__nand2_1 _4333_ (.A(_0185_),
    .B(_0253_),
    .Y(_0254_));
 sky130_fd_sc_hs__o211ai_2 _4334_ (.A1(_0181_),
    .A2(_0185_),
    .B1(_0252_),
    .C1(_0254_),
    .Y(_0255_));
 sky130_fd_sc_hs__a311oi_4 _4335_ (.A1(_0181_),
    .A2(_0180_),
    .A3(_0185_),
    .B1(_0250_),
    .C1(_0255_),
    .Y(net14));
 sky130_fd_sc_hs__inv_1 _4336_ (.A(_0192_),
    .Y(_0256_));
 sky130_fd_sc_hs__nand3_1 _4337_ (.A(_0192_),
    .B(_0124_),
    .C(_0130_),
    .Y(_0257_));
 sky130_fd_sc_hs__a211oi_4 _4338_ (.A1(_0164_),
    .A2(_0173_),
    .B1(_0179_),
    .C1(_0257_),
    .Y(_0258_));
 sky130_fd_sc_hs__nor2_1 _4339_ (.A(_0192_),
    .B(_0130_),
    .Y(_0259_));
 sky130_fd_sc_hs__o211ai_1 _4340_ (.A1(_0129_),
    .A2(_0187_),
    .B1(_0188_),
    .C1(_0259_),
    .Y(_0260_));
 sky130_fd_sc_hs__nor2_1 _4341_ (.A(_0192_),
    .B(_0124_),
    .Y(_0261_));
 sky130_fd_sc_hs__o211ai_1 _4342_ (.A1(_0129_),
    .A2(_0187_),
    .B1(_0188_),
    .C1(_0261_),
    .Y(_0262_));
 sky130_fd_sc_hs__o211ai_1 _4343_ (.A1(_0256_),
    .A2(_0189_),
    .B1(_0260_),
    .C1(_0262_),
    .Y(_0263_));
 sky130_fd_sc_hs__a311oi_4 _4344_ (.A1(_0256_),
    .A2(_0180_),
    .A3(_0189_),
    .B1(_0258_),
    .C1(_0263_),
    .Y(net211));
 sky130_fd_sc_hs__or4_2 _4345_ (.A(net209),
    .B(net208),
    .C(net207),
    .D(net211),
    .X(_0264_));
 sky130_fd_sc_hs__a31o_4 _4346_ (.A1(_0233_),
    .A2(_0240_),
    .A3(_0242_),
    .B1(_0160_),
    .X(_0265_));
 sky130_fd_sc_hs__a21oi_2 _4347_ (.A1(_3673_),
    .A2(_3668_),
    .B1(_3672_),
    .Y(_0266_));
 sky130_fd_sc_hs__nand2_1 _4348_ (.A(_3677_),
    .B(_0128_),
    .Y(_0267_));
 sky130_fd_sc_hs__a21oi_1 _4349_ (.A1(_0128_),
    .A2(_3676_),
    .B1(_3680_),
    .Y(_0268_));
 sky130_fd_sc_hs__o21ai_2 _4350_ (.A1(_0266_),
    .A2(_0267_),
    .B1(_0268_),
    .Y(_0269_));
 sky130_fd_sc_hs__or3b_4 _4351_ (.A(_0218_),
    .B(_0269_),
    .C_N(_0230_),
    .X(_0270_));
 sky130_fd_sc_hs__or3b_1 _4352_ (.A(_3684_),
    .B(_3688_),
    .C_N(_3693_),
    .X(_0271_));
 sky130_fd_sc_hs__a21oi_1 _4353_ (.A1(_0125_),
    .A2(_0266_),
    .B1(_0182_),
    .Y(_0272_));
 sky130_fd_sc_hs__o21a_1 _4354_ (.A1(_3676_),
    .A2(_0272_),
    .B1(_0128_),
    .X(_0273_));
 sky130_fd_sc_hs__nor3_4 _4355_ (.A(_0218_),
    .B(_0234_),
    .C(_0269_),
    .Y(_0274_));
 sky130_fd_sc_hs__a2bb2oi_4 _4356_ (.A1_N(_3680_),
    .A2_N(_0273_),
    .B1(_0274_),
    .B2(_0230_),
    .Y(_0275_));
 sky130_fd_sc_hs__o21ai_1 _4357_ (.A1(_3685_),
    .A2(_3684_),
    .B1(_0192_),
    .Y(_0276_));
 sky130_fd_sc_hs__nand3b_1 _4358_ (.A_N(_3688_),
    .B(_0276_),
    .C(_3693_),
    .Y(_0277_));
 sky130_fd_sc_hs__nand3b_1 _4359_ (.A_N(_3693_),
    .B(_3684_),
    .C(_0192_),
    .Y(_0278_));
 sky130_fd_sc_hs__nand2b_1 _4360_ (.A_N(_3693_),
    .B(_3688_),
    .Y(_0279_));
 sky130_fd_sc_hs__o2111a_1 _4361_ (.A1(_0275_),
    .A2(_0271_),
    .B1(_0277_),
    .C1(_0278_),
    .D1(_0279_),
    .X(_0280_));
 sky130_fd_sc_hs__nor2_1 _4362_ (.A(_3693_),
    .B(_0276_),
    .Y(_0281_));
 sky130_fd_sc_hs__o211ai_1 _4363_ (.A1(_0265_),
    .A2(_0270_),
    .B1(_0281_),
    .C1(_0275_),
    .Y(_0282_));
 sky130_fd_sc_hs__o311ai_2 _4364_ (.A1(_0265_),
    .A2(_0270_),
    .A3(_0271_),
    .B1(_0280_),
    .C1(_0282_),
    .Y(net10));
 sky130_fd_sc_hs__xor2_4 _4365_ (.A(_0126_),
    .B(_0211_),
    .X(net205));
 sky130_fd_sc_hs__nor4b_4 _4366_ (.A(_3600_),
    .B(_0236_),
    .C(_0237_),
    .D_N(_0238_),
    .Y(_0283_));
 sky130_fd_sc_hs__nand2_1 _4367_ (.A(_0238_),
    .B(_0241_),
    .Y(_0284_));
 sky130_fd_sc_hs__a21oi_4 _4368_ (.A1(_0200_),
    .A2(_0238_),
    .B1(_0155_),
    .Y(_0285_));
 sky130_fd_sc_hs__nand2_2 _4369_ (.A(_0284_),
    .B(_0285_),
    .Y(_0286_));
 sky130_fd_sc_hs__nand3_2 _4370_ (.A(_0154_),
    .B(_3621_),
    .C(_3612_),
    .Y(_0287_));
 sky130_fd_sc_hs__a21oi_2 _4371_ (.A1(_3621_),
    .A2(_3616_),
    .B1(_3620_),
    .Y(_0288_));
 sky130_fd_sc_hs__nand2_4 _4372_ (.A(_0287_),
    .B(_0288_),
    .Y(_0289_));
 sky130_fd_sc_hs__a21oi_4 _4373_ (.A1(_0163_),
    .A2(_0289_),
    .B1(_0166_),
    .Y(_0290_));
 sky130_fd_sc_hs__inv_2 _4374_ (.A(_0177_),
    .Y(_0291_));
 sky130_fd_sc_hs__o211a_1 _4375_ (.A1(_0283_),
    .A2(_0286_),
    .B1(_0290_),
    .C1(_0291_),
    .X(_0292_));
 sky130_fd_sc_hs__or3_1 _4376_ (.A(_0177_),
    .B(_0163_),
    .C(_0166_),
    .X(_0293_));
 sky130_fd_sc_hs__o21ai_2 _4377_ (.A1(_0291_),
    .A2(_0290_),
    .B1(_0293_),
    .Y(_0294_));
 sky130_fd_sc_hs__nor4_4 _4378_ (.A(_0291_),
    .B(_0153_),
    .C(_0283_),
    .D(_0286_),
    .Y(_0295_));
 sky130_fd_sc_hs__nor3_4 _4379_ (.A(_0292_),
    .B(_0294_),
    .C(_0295_),
    .Y(net15));
 sky130_fd_sc_hs__nor3b_1 _4380_ (.A(_0169_),
    .B(_0207_),
    .C_N(_0203_),
    .Y(_0296_));
 sky130_fd_sc_hs__and3_1 _4381_ (.A(_3613_),
    .B(_0240_),
    .C(_0242_),
    .X(_0297_));
 sky130_fd_sc_hs__a21oi_2 _4382_ (.A1(_0240_),
    .A2(_0242_),
    .B1(_3613_),
    .Y(_0298_));
 sky130_fd_sc_hs__or2_4 _4383_ (.A(_0297_),
    .B(_0298_),
    .X(_0299_));
 sky130_fd_sc_hs__clkinv_8 _4384_ (.A(_0299_),
    .Y(net222));
 sky130_fd_sc_hs__or2_2 _4385_ (.A(_0236_),
    .B(_0237_),
    .X(_0300_));
 sky130_fd_sc_hs__a21oi_4 _4386_ (.A1(_3601_),
    .A2(_0300_),
    .B1(_3600_),
    .Y(_0301_));
 sky130_fd_sc_hs__xnor2_4 _4387_ (.A(_3605_),
    .B(_0301_),
    .Y(net220));
 sky130_fd_sc_hs__and2_2 _4388_ (.A(_0143_),
    .B(_0144_),
    .X(_0302_));
 sky130_fd_sc_hs__a22oi_4 _4389_ (.A1(_0137_),
    .A2(_0138_),
    .B1(_0136_),
    .B2(_0302_),
    .Y(_0303_));
 sky130_fd_sc_hs__xor2_4 _4390_ (.A(_3593_),
    .B(_0303_),
    .X(net217));
 sky130_fd_sc_hs__nand2_1 _4391_ (.A(_0168_),
    .B(_0204_),
    .Y(_0304_));
 sky130_fd_sc_hs__mux2i_4 _4392_ (.A0(_0304_),
    .A1(_0168_),
    .S(_0207_),
    .Y(_0305_));
 sky130_fd_sc_hs__xnor2_4 _4393_ (.A(_3581_),
    .B(_2229_),
    .Y(_0306_));
 sky130_fd_sc_hs__clkinv_8 _4394_ (.A(_0306_),
    .Y(net202));
 sky130_fd_sc_hs__a21o_1 _4395_ (.A1(_3581_),
    .A2(_2229_),
    .B1(_3580_),
    .X(_0307_));
 sky130_fd_sc_hs__a21oi_4 _4396_ (.A1(_3585_),
    .A2(_0307_),
    .B1(_3584_),
    .Y(_0308_));
 sky130_fd_sc_hs__xnor2_4 _4397_ (.A(_3589_),
    .B(_0308_),
    .Y(net216));
 sky130_fd_sc_hs__nor4_4 _4398_ (.A(net191),
    .B(_0305_),
    .C(net202),
    .D(net216),
    .Y(_0309_));
 sky130_fd_sc_hs__nand4_2 _4399_ (.A(_0117_),
    .B(_0119_),
    .C(_0120_),
    .D(_0135_),
    .Y(_0310_));
 sky130_fd_sc_hs__o211ai_4 _4400_ (.A1(_0111_),
    .A2(_0113_),
    .B1(_0135_),
    .C1(_0115_),
    .Y(_0311_));
 sky130_fd_sc_hs__nand2_1 _4401_ (.A(_0132_),
    .B(_0135_),
    .Y(_0312_));
 sky130_fd_sc_hs__nand4_2 _4402_ (.A(_0310_),
    .B(_0311_),
    .C(_0312_),
    .D(_0143_),
    .Y(_0313_));
 sky130_fd_sc_hs__xnor2_4 _4403_ (.A(_3585_),
    .B(_0313_),
    .Y(_0314_));
 sky130_fd_sc_hs__o21ai_1 _4404_ (.A1(_0138_),
    .A2(_0235_),
    .B1(_0137_),
    .Y(_0315_));
 sky130_fd_sc_hs__a21oi_4 _4405_ (.A1(_3593_),
    .A2(_0315_),
    .B1(_3592_),
    .Y(_0316_));
 sky130_fd_sc_hs__xor2_4 _4406_ (.A(_3597_),
    .B(_0316_),
    .X(_0317_));
 sky130_fd_sc_hs__nand3_1 _4407_ (.A(_0309_),
    .B(_0314_),
    .C(_0317_),
    .Y(_0318_));
 sky130_fd_sc_hs__or4_1 _4408_ (.A(net222),
    .B(net220),
    .C(net217),
    .D(_0318_),
    .X(_0319_));
 sky130_fd_sc_hs__nor3_1 _4409_ (.A(net197),
    .B(_0296_),
    .C(_0319_),
    .Y(_0320_));
 sky130_fd_sc_hs__nand4_2 _4410_ (.A(_0310_),
    .B(_0311_),
    .C(_0312_),
    .D(_0302_),
    .Y(_0321_));
 sky130_fd_sc_hs__a21oi_1 _4411_ (.A1(_0140_),
    .A2(_0321_),
    .B1(_0142_),
    .Y(_0322_));
 sky130_fd_sc_hs__nand2_1 _4412_ (.A(_3601_),
    .B(_0148_),
    .Y(_0323_));
 sky130_fd_sc_hs__o21ai_1 _4413_ (.A1(_0322_),
    .A2(_0323_),
    .B1(_0159_),
    .Y(_0324_));
 sky130_fd_sc_hs__nor2_1 _4414_ (.A(_0149_),
    .B(_0165_),
    .Y(_0325_));
 sky130_fd_sc_hs__o2111a_1 _4415_ (.A1(_0322_),
    .A2(_0323_),
    .B1(_0325_),
    .C1(_0159_),
    .D1(_0161_),
    .X(_0326_));
 sky130_fd_sc_hs__nand2_1 _4416_ (.A(_3625_),
    .B(_3629_),
    .Y(_0327_));
 sky130_fd_sc_hs__a21oi_1 _4417_ (.A1(_0161_),
    .A2(_0155_),
    .B1(_0327_),
    .Y(_0328_));
 sky130_fd_sc_hs__nor2_1 _4418_ (.A(_0327_),
    .B(_0161_),
    .Y(_0329_));
 sky130_fd_sc_hs__o21ai_1 _4419_ (.A1(_0165_),
    .A2(_0329_),
    .B1(_0149_),
    .Y(_0330_));
 sky130_fd_sc_hs__o31ai_1 _4420_ (.A1(_0149_),
    .A2(_0165_),
    .A3(_0328_),
    .B1(_0330_),
    .Y(_0331_));
 sky130_fd_sc_hs__a211oi_4 _4421_ (.A1(_0156_),
    .A2(_0324_),
    .B1(_0326_),
    .C1(_0331_),
    .Y(net16));
 sky130_fd_sc_hs__o211ai_4 _4422_ (.A1(_0136_),
    .A2(_0141_),
    .B1(_0146_),
    .C1(_0159_),
    .Y(_0332_));
 sky130_fd_sc_hs__a211oi_4 _4423_ (.A1(_0285_),
    .A2(_0332_),
    .B1(_3625_),
    .C1(_0289_),
    .Y(_0333_));
 sky130_fd_sc_hs__nor3_1 _4424_ (.A(_0150_),
    .B(_0155_),
    .C(_0200_),
    .Y(_0334_));
 sky130_fd_sc_hs__a22o_4 _4425_ (.A1(_3625_),
    .A2(_0162_),
    .B1(_0147_),
    .B2(_0334_),
    .X(_0335_));
 sky130_fd_sc_hs__nor2_8 _4426_ (.A(_0333_),
    .B(_0335_),
    .Y(net194));
 sky130_fd_sc_hs__a211oi_4 _4427_ (.A1(_0140_),
    .A2(_0321_),
    .B1(_3601_),
    .C1(_0142_),
    .Y(_0336_));
 sky130_fd_sc_hs__nor2_8 _4428_ (.A(_0147_),
    .B(_0336_),
    .Y(net219));
 sky130_fd_sc_hs__o21bai_1 _4429_ (.A1(_0157_),
    .A2(_0158_),
    .B1_N(_3608_),
    .Y(_0337_));
 sky130_fd_sc_hs__nor3b_2 _4430_ (.A(_3612_),
    .B(_0337_),
    .C_N(_0154_),
    .Y(_0338_));
 sky130_fd_sc_hs__clkinv_2 _4431_ (.A(_3613_),
    .Y(_0339_));
 sky130_fd_sc_hs__nor3_4 _4432_ (.A(_0339_),
    .B(_0154_),
    .C(_0200_),
    .Y(_0340_));
 sky130_fd_sc_hs__mux2i_4 _4433_ (.A0(_0338_),
    .A1(_0340_),
    .S(_0147_),
    .Y(_0341_));
 sky130_fd_sc_hs__nor2_2 _4434_ (.A(_0339_),
    .B(_0159_),
    .Y(_0342_));
 sky130_fd_sc_hs__a21oi_1 _4435_ (.A1(_0200_),
    .A2(_0238_),
    .B1(_0339_),
    .Y(_0343_));
 sky130_fd_sc_hs__o21ai_1 _4436_ (.A1(_3612_),
    .A2(_0343_),
    .B1(_0154_),
    .Y(_0344_));
 sky130_fd_sc_hs__o31ai_4 _4437_ (.A1(_0154_),
    .A2(_3612_),
    .A3(_0342_),
    .B1(_0344_),
    .Y(_0345_));
 sky130_fd_sc_hs__nand2_8 _4438_ (.A(_0341_),
    .B(_0345_),
    .Y(net192));
 sky130_fd_sc_hs__nor4_2 _4439_ (.A(net196),
    .B(net194),
    .C(net219),
    .D(net192),
    .Y(_0346_));
 sky130_fd_sc_hs__nor2_1 _4440_ (.A(_3605_),
    .B(_3604_),
    .Y(_0347_));
 sky130_fd_sc_hs__nor3_2 _4441_ (.A(_3601_),
    .B(_3600_),
    .C(_3604_),
    .Y(_0348_));
 sky130_fd_sc_hs__a2111oi_4 _4442_ (.A1(_0140_),
    .A2(_0321_),
    .B1(_3600_),
    .C1(_3604_),
    .D1(_0142_),
    .Y(_0349_));
 sky130_fd_sc_hs__or4_1 _4443_ (.A(_0157_),
    .B(_0347_),
    .C(_0348_),
    .D(_0349_),
    .X(_0350_));
 sky130_fd_sc_hs__o31ai_2 _4444_ (.A1(_0347_),
    .A2(_0348_),
    .A3(_0349_),
    .B1(_0157_),
    .Y(_0351_));
 sky130_fd_sc_hs__and2_4 _4445_ (.A(_0350_),
    .B(_0351_),
    .X(net221));
 sky130_fd_sc_hs__nor3_1 _4446_ (.A(_0168_),
    .B(_0203_),
    .C(_0204_),
    .Y(_0352_));
 sky130_fd_sc_hs__nor2_1 _4447_ (.A(net221),
    .B(_0352_),
    .Y(_0353_));
 sky130_fd_sc_hs__nand4b_1 _4448_ (.A_N(net205),
    .B(_0320_),
    .C(_0346_),
    .D(_0353_),
    .Y(_0354_));
 sky130_fd_sc_hs__o21bai_1 _4449_ (.A1(_0174_),
    .A2(_0222_),
    .B1_N(_3652_),
    .Y(_0355_));
 sky130_fd_sc_hs__nand2_1 _4450_ (.A(_0177_),
    .B(_0175_),
    .Y(_0356_));
 sky130_fd_sc_hs__and2_1 _4451_ (.A(_0284_),
    .B(_0285_),
    .X(_0357_));
 sky130_fd_sc_hs__nand2_1 _4452_ (.A(_0240_),
    .B(_0357_),
    .Y(_0358_));
 sky130_fd_sc_hs__o21a_1 _4453_ (.A1(_0356_),
    .A2(_0290_),
    .B1(_0220_),
    .X(_0359_));
 sky130_fd_sc_hs__o31ai_4 _4454_ (.A1(_0153_),
    .A2(_0356_),
    .A3(_0358_),
    .B1(_0359_),
    .Y(_0360_));
 sky130_fd_sc_hs__nand2_1 _4455_ (.A(_0167_),
    .B(_3657_),
    .Y(_0361_));
 sky130_fd_sc_hs__nor2_2 _4456_ (.A(_0221_),
    .B(_0361_),
    .Y(_0362_));
 sky130_fd_sc_hs__a221oi_4 _4457_ (.A1(_3657_),
    .A2(_0355_),
    .B1(_0360_),
    .B2(_0362_),
    .C1(_3656_),
    .Y(_0363_));
 sky130_fd_sc_hs__xnor2_4 _4458_ (.A(_3661_),
    .B(_0363_),
    .Y(net204));
 sky130_fd_sc_hs__xor2_4 _4459_ (.A(_3645_),
    .B(_0360_),
    .X(net199));
 sky130_fd_sc_hs__xnor2_4 _4460_ (.A(_3657_),
    .B(_0180_),
    .Y(net203));
 sky130_fd_sc_hs__a21oi_4 _4461_ (.A1(_0149_),
    .A2(_0165_),
    .B1(_3632_),
    .Y(_0364_));
 sky130_fd_sc_hs__a211o_1 _4462_ (.A1(_0164_),
    .A2(_0364_),
    .B1(_0291_),
    .C1(_0175_),
    .X(_0365_));
 sky130_fd_sc_hs__nand4b_2 _4463_ (.A_N(_3636_),
    .B(_0164_),
    .C(_0364_),
    .D(_0175_),
    .Y(_0366_));
 sky130_fd_sc_hs__inv_1 _4464_ (.A(_0175_),
    .Y(_0367_));
 sky130_fd_sc_hs__nor3_2 _4465_ (.A(_0177_),
    .B(_0367_),
    .C(_3636_),
    .Y(_0368_));
 sky130_fd_sc_hs__a21oi_4 _4466_ (.A1(_0367_),
    .A2(_3636_),
    .B1(_0368_),
    .Y(_0369_));
 sky130_fd_sc_hs__a21oi_1 _4467_ (.A1(_0240_),
    .A2(_0357_),
    .B1(_0289_),
    .Y(_0370_));
 sky130_fd_sc_hs__a2111o_1 _4468_ (.A1(_0240_),
    .A2(_0357_),
    .B1(_0151_),
    .C1(_3624_),
    .D1(_0289_),
    .X(_0371_));
 sky130_fd_sc_hs__nor3_1 _4469_ (.A(_3625_),
    .B(_0151_),
    .C(_3624_),
    .Y(_0372_));
 sky130_fd_sc_hs__a21oi_1 _4470_ (.A1(_0151_),
    .A2(_3624_),
    .B1(_0372_),
    .Y(_0373_));
 sky130_fd_sc_hs__o311a_4 _4471_ (.A1(_0150_),
    .A2(_3629_),
    .A3(_0370_),
    .B1(_0371_),
    .C1(_0373_),
    .X(_0374_));
 sky130_fd_sc_hs__nand4_2 _4472_ (.A(_0365_),
    .B(_0366_),
    .C(_0369_),
    .D(_0374_),
    .Y(_0375_));
 sky130_fd_sc_hs__nor4_4 _4473_ (.A(net204),
    .B(net199),
    .C(net203),
    .D(_0375_),
    .Y(_0376_));
 sky130_fd_sc_hs__o21ai_4 _4474_ (.A1(_0265_),
    .A2(_0270_),
    .B1(_0275_),
    .Y(_0377_));
 sky130_fd_sc_hs__buf_8 _4475_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .X(_0378_));
 sky130_fd_sc_hs__nor4_4 _4476_ (.A(_0102_),
    .B(\genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .C(_0378_),
    .D(\genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .Y(_0379_));
 sky130_fd_sc_hs__nor2b_2 _4477_ (.A(net177),
    .B_N(net366),
    .Y(_0380_));
 sky130_fd_sc_hs__clkinv_8 _4478_ (.A(_0378_),
    .Y(_0381_));
 sky130_fd_sc_hs__buf_8 _4479_ (.A(net113),
    .X(_0382_));
 sky130_fd_sc_hs__inv_8 _4480_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .Y(_0383_));
 sky130_fd_sc_hs__o22ai_4 _4481_ (.A1(_0381_),
    .A2(_0382_),
    .B1(net145),
    .B2(_0383_),
    .Y(_0384_));
 sky130_fd_sc_hs__inv_2 _4482_ (.A(net113),
    .Y(_0385_));
 sky130_fd_sc_hs__clkbuf_16 _4483_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .X(_0386_));
 sky130_fd_sc_hs__nor2_8 _4484_ (.A(_0102_),
    .B(_0386_),
    .Y(_0387_));
 sky130_fd_sc_hs__a21oi_1 _4485_ (.A1(_0385_),
    .A2(net105),
    .B1(_0387_),
    .Y(_0388_));
 sky130_fd_sc_hs__nor3_1 _4486_ (.A(_0380_),
    .B(_0384_),
    .C(_0388_),
    .Y(_0389_));
 sky130_fd_sc_hs__inv_1 _4487_ (.A(net105),
    .Y(_0390_));
 sky130_fd_sc_hs__clkinv_8 _4488_ (.A(_0102_),
    .Y(_0391_));
 sky130_fd_sc_hs__clkinv_8 _4489_ (.A(_0386_),
    .Y(_0392_));
 sky130_fd_sc_hs__nand2_4 _4490_ (.A(_0391_),
    .B(_0392_),
    .Y(_0393_));
 sky130_fd_sc_hs__o211a_1 _4491_ (.A1(_0390_),
    .A2(_0384_),
    .B1(_0393_),
    .C1(_0382_),
    .X(_0394_));
 sky130_fd_sc_hs__o21a_1 _4492_ (.A1(_0389_),
    .A2(_0394_),
    .B1(_0132_),
    .X(_0395_));
 sky130_fd_sc_hs__xnor2_4 _4493_ (.A(net66),
    .B(net34),
    .Y(_0396_));
 sky130_fd_sc_hs__nor3_4 _4494_ (.A(_0133_),
    .B(_0134_),
    .C(_0396_),
    .Y(_0397_));
 sky130_fd_sc_hs__o21ai_1 _4495_ (.A1(_0133_),
    .A2(_0134_),
    .B1(_0396_),
    .Y(_0398_));
 sky130_fd_sc_hs__nor3b_4 _4496_ (.A(_0132_),
    .B(_0397_),
    .C_N(_0398_),
    .Y(_0399_));
 sky130_fd_sc_hs__nor2_4 _4497_ (.A(_0395_),
    .B(_0399_),
    .Y(_0400_));
 sky130_fd_sc_hs__nand2_1 _4498_ (.A(_0192_),
    .B(_3684_),
    .Y(_0401_));
 sky130_fd_sc_hs__a211oi_2 _4499_ (.A1(_3697_),
    .A2(_3692_),
    .B1(_3696_),
    .C1(_3688_),
    .Y(_0402_));
 sky130_fd_sc_hs__and2_1 _4500_ (.A(_0401_),
    .B(_0402_),
    .X(_0403_));
 sky130_fd_sc_hs__and3_2 _4501_ (.A(_0377_),
    .B(_0400_),
    .C(_0403_),
    .X(_0404_));
 sky130_fd_sc_hs__nand2b_1 _4502_ (.A_N(_3688_),
    .B(_0276_),
    .Y(_0405_));
 sky130_fd_sc_hs__a21o_1 _4503_ (.A1(_3693_),
    .A2(_0405_),
    .B1(_3692_),
    .X(_0406_));
 sky130_fd_sc_hs__a21oi_4 _4504_ (.A1(_3697_),
    .A2(_0406_),
    .B1(_3696_),
    .Y(_0407_));
 sky130_fd_sc_hs__and2_2 _4505_ (.A(_0400_),
    .B(_0407_),
    .X(_0408_));
 sky130_fd_sc_hs__a211oi_4 _4506_ (.A1(_0377_),
    .A2(_0403_),
    .B1(_0407_),
    .C1(_0400_),
    .Y(_0409_));
 sky130_fd_sc_hs__or3_1 _4507_ (.A(_0404_),
    .B(_0408_),
    .C(_0409_),
    .X(_0410_));
 sky130_fd_sc_hs__clkbuf_16 _4508_ (.A(_0410_),
    .X(net215));
 sky130_fd_sc_hs__nor2_1 _4509_ (.A(_0283_),
    .B(_0286_),
    .Y(_0411_));
 sky130_fd_sc_hs__nand3b_1 _4510_ (.A_N(_0223_),
    .B(_0290_),
    .C(_0174_),
    .Y(_0412_));
 sky130_fd_sc_hs__nor3_1 _4511_ (.A(_0167_),
    .B(_0223_),
    .C(_0228_),
    .Y(_0413_));
 sky130_fd_sc_hs__nor4_2 _4512_ (.A(_0167_),
    .B(_0163_),
    .C(_0166_),
    .D(_0223_),
    .Y(_0414_));
 sky130_fd_sc_hs__a211oi_1 _4513_ (.A1(_0167_),
    .A2(_0223_),
    .B1(_0413_),
    .C1(_0414_),
    .Y(_0415_));
 sky130_fd_sc_hs__and3_1 _4514_ (.A(_0167_),
    .B(_0163_),
    .C(_0228_),
    .X(_0416_));
 sky130_fd_sc_hs__a21bo_1 _4515_ (.A1(_0287_),
    .A2(_0288_),
    .B1_N(_0163_),
    .X(_0417_));
 sky130_fd_sc_hs__nand2_1 _4516_ (.A(_0167_),
    .B(_0228_),
    .Y(_0418_));
 sky130_fd_sc_hs__a21oi_1 _4517_ (.A1(_0417_),
    .A2(_0364_),
    .B1(_0418_),
    .Y(_0419_));
 sky130_fd_sc_hs__a31oi_1 _4518_ (.A1(_0240_),
    .A2(_0357_),
    .A3(_0416_),
    .B1(_0419_),
    .Y(_0420_));
 sky130_fd_sc_hs__o211a_2 _4519_ (.A1(_0411_),
    .A2(_0412_),
    .B1(_0415_),
    .C1(_0420_),
    .X(_0421_));
 sky130_fd_sc_hs__buf_16 _4520_ (.A(_0421_),
    .X(net201));
 sky130_fd_sc_hs__nand3_4 _4521_ (.A(_0231_),
    .B(_0243_),
    .C(_0245_),
    .Y(_0422_));
 sky130_fd_sc_hs__xor2_4 _4522_ (.A(_3669_),
    .B(_0422_),
    .X(net206));
 sky130_fd_sc_hs__xor2_4 _4523_ (.A(_3621_),
    .B(_0265_),
    .X(net193));
 sky130_fd_sc_hs__xnor2_4 _4524_ (.A(_3685_),
    .B(_0377_),
    .Y(net210));
 sky130_fd_sc_hs__or4_1 _4525_ (.A(net201),
    .B(net206),
    .C(net365),
    .D(net210),
    .X(_0423_));
 sky130_fd_sc_hs__nor2_2 _4526_ (.A(net215),
    .B(_0423_),
    .Y(_0424_));
 sky130_fd_sc_hs__nand4bb_4 _4527_ (.A_N(net11),
    .B_N(_0354_),
    .C(_0376_),
    .D(_0424_),
    .Y(_0425_));
 sky130_fd_sc_hs__or4_4 _4528_ (.A(net78),
    .B(net214),
    .C(_0264_),
    .D(_0425_),
    .X(_0426_));
 sky130_fd_sc_hs__clkbuf_16 _4529_ (.A(_0383_),
    .X(_0427_));
 sky130_fd_sc_hs__nor2_1 _4530_ (.A(_0427_),
    .B(_0094_),
    .Y(_0428_));
 sky130_fd_sc_hs__a31o_1 _4531_ (.A1(_0123_),
    .A2(_0094_),
    .A3(_0426_),
    .B1(_0428_),
    .X(_0004_));
 sky130_fd_sc_hs__nand2_1 _4532_ (.A(_0123_),
    .B(net79),
    .Y(_0429_));
 sky130_fd_sc_hs__buf_8 _4533_ (.A(_0378_),
    .X(_0430_));
 sky130_fd_sc_hs__a21oi_1 _4534_ (.A1(net187),
    .A2(net79),
    .B1(_0092_),
    .Y(_0431_));
 sky130_fd_sc_hs__a21oi_1 _4535_ (.A1(_0430_),
    .A2(net79),
    .B1(_0431_),
    .Y(_0432_));
 sky130_fd_sc_hs__o21ai_1 _4536_ (.A1(_0426_),
    .A2(_0429_),
    .B1(_0432_),
    .Y(_0003_));
 sky130_fd_sc_hs__buf_8 _4537_ (.A(_0391_),
    .X(_0433_));
 sky130_fd_sc_hs__o22ai_1 _4538_ (.A1(_0392_),
    .A2(_0094_),
    .B1(_0101_),
    .B2(_0433_),
    .Y(_0002_));
 sky130_fd_sc_hs__a21oi_1 _4539_ (.A1(net187),
    .A2(net120),
    .B1(\genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0] ),
    .Y(_0434_));
 sky130_fd_sc_hs__a21oi_1 _4540_ (.A1(net120),
    .A2(_0087_),
    .B1(_0434_),
    .Y(_0000_));
 sky130_fd_sc_hs__clkbuf_16 _4541_ (.A(imd_val_q_i[34]),
    .X(_0435_));
 sky130_fd_sc_hs__buf_8 _4542_ (.A(imd_val_q_i[50]),
    .X(_0436_));
 sky130_fd_sc_hs__mux2_1 _4543_ (.A0(_0435_),
    .A1(_0436_),
    .S(_0083_),
    .X(_0437_));
 sky130_fd_sc_hs__or2_4 _4544_ (.A(_0081_),
    .B(\genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[2] ),
    .X(_0438_));
 sky130_fd_sc_hs__buf_16 _4545_ (.A(_0438_),
    .X(_0439_));
 sky130_fd_sc_hs__clkbuf_16 _4546_ (.A(_0439_),
    .X(_0440_));
 sky130_fd_sc_hs__a22o_1 _4547_ (.A1(_0084_),
    .A2(_0437_),
    .B1(_0440_),
    .B2(_0436_),
    .X(_3699_));
 sky130_fd_sc_hs__mux2i_4 _4548_ (.A0(net153),
    .A1(net160),
    .S(_0438_),
    .Y(_0441_));
 sky130_fd_sc_hs__clkbuf_8 _4549_ (.A(_0441_),
    .X(_0442_));
 sky130_fd_sc_hs__nor2_8 _4550_ (.A(_0081_),
    .B(_0084_),
    .Y(_0443_));
 sky130_fd_sc_hs__mux2i_4 _4551_ (.A0(net128),
    .A1(net121),
    .S(_0443_),
    .Y(_0444_));
 sky130_fd_sc_hs__buf_8 _4552_ (.A(_0444_),
    .X(_0445_));
 sky130_fd_sc_hs__nor2_2 _4553_ (.A(_0442_),
    .B(_0445_),
    .Y(_3698_));
 sky130_fd_sc_hs__buf_8 _4554_ (.A(imd_val_q_i[51]),
    .X(_0446_));
 sky130_fd_sc_hs__buf_8 _4555_ (.A(imd_val_q_i[35]),
    .X(_0447_));
 sky130_fd_sc_hs__mux2_1 _4556_ (.A0(_0447_),
    .A1(_0446_),
    .S(_0083_),
    .X(_0448_));
 sky130_fd_sc_hs__a22oi_4 _4557_ (.A1(_0446_),
    .A2(_0440_),
    .B1(_0448_),
    .B2(_0084_),
    .Y(_2232_));
 sky130_fd_sc_hs__buf_8 _4558_ (.A(imd_val_q_i[52]),
    .X(_0449_));
 sky130_fd_sc_hs__clkbuf_16 _4559_ (.A(imd_val_q_i[36]),
    .X(_0450_));
 sky130_fd_sc_hs__mux2_1 _4560_ (.A0(_0450_),
    .A1(_0449_),
    .S(_0083_),
    .X(_0451_));
 sky130_fd_sc_hs__a22oi_4 _4561_ (.A1(_0449_),
    .A2(_0440_),
    .B1(_0451_),
    .B2(_0084_),
    .Y(_2237_));
 sky130_fd_sc_hs__mux2i_4 _4562_ (.A0(net175),
    .A1(net162),
    .S(_0439_),
    .Y(_0452_));
 sky130_fd_sc_hs__buf_4 _4563_ (.A(_0452_),
    .X(_0453_));
 sky130_fd_sc_hs__nor2_2 _4564_ (.A(_0445_),
    .B(_0453_),
    .Y(_2240_));
 sky130_fd_sc_hs__buf_16 _4565_ (.A(_0443_),
    .X(_0454_));
 sky130_fd_sc_hs__mux2i_4 _4566_ (.A0(net131),
    .A1(net146),
    .S(_0454_),
    .Y(_0455_));
 sky130_fd_sc_hs__clkbuf_8 _4567_ (.A(_0455_),
    .X(_0456_));
 sky130_fd_sc_hs__nor2_2 _4568_ (.A(_0442_),
    .B(_0456_),
    .Y(_2246_));
 sky130_fd_sc_hs__mux2i_4 _4569_ (.A0(net130),
    .A1(net143),
    .S(_0454_),
    .Y(_0457_));
 sky130_fd_sc_hs__clkbuf_8 _4570_ (.A(_0457_),
    .X(_0458_));
 sky130_fd_sc_hs__mux2i_4 _4571_ (.A0(net164),
    .A1(net161),
    .S(_0439_),
    .Y(_0459_));
 sky130_fd_sc_hs__clkbuf_8 _4572_ (.A(_0459_),
    .X(_0460_));
 sky130_fd_sc_hs__nor2_1 _4573_ (.A(_0458_),
    .B(_0460_),
    .Y(_2245_));
 sky130_fd_sc_hs__mux2i_4 _4574_ (.A0(net129),
    .A1(net132),
    .S(_0454_),
    .Y(_0461_));
 sky130_fd_sc_hs__clkbuf_8 _4575_ (.A(_0461_),
    .X(_0462_));
 sky130_fd_sc_hs__nor2_1 _4576_ (.A(_0453_),
    .B(_0462_),
    .Y(_3720_));
 sky130_fd_sc_hs__mux2i_4 _4577_ (.A0(net178),
    .A1(net163),
    .S(_0439_),
    .Y(_0463_));
 sky130_fd_sc_hs__buf_4 _4578_ (.A(_0463_),
    .X(_0464_));
 sky130_fd_sc_hs__nor2_1 _4579_ (.A(_0445_),
    .B(_0464_),
    .Y(_3719_));
 sky130_fd_sc_hs__mux2i_4 _4580_ (.A0(net133),
    .A1(net147),
    .S(_0443_),
    .Y(_0465_));
 sky130_fd_sc_hs__clkbuf_8 _4581_ (.A(_0465_),
    .X(_0466_));
 sky130_fd_sc_hs__nor2_2 _4582_ (.A(_0442_),
    .B(_0466_),
    .Y(_2255_));
 sky130_fd_sc_hs__nor2_2 _4583_ (.A(_0456_),
    .B(_0460_),
    .Y(_2254_));
 sky130_fd_sc_hs__nor2_1 _4584_ (.A(_0453_),
    .B(_0458_),
    .Y(_2261_));
 sky130_fd_sc_hs__nor2_1 _4585_ (.A(_0462_),
    .B(_0464_),
    .Y(_2260_));
 sky130_fd_sc_hs__mux2i_4 _4586_ (.A0(net179),
    .A1(net165),
    .S(_0439_),
    .Y(_0467_));
 sky130_fd_sc_hs__clkbuf_8 _4587_ (.A(_0467_),
    .X(_0468_));
 sky130_fd_sc_hs__nor2_1 _4588_ (.A(_0445_),
    .B(_0468_),
    .Y(_2259_));
 sky130_fd_sc_hs__mux2i_4 _4589_ (.A0(net134),
    .A1(net148),
    .S(_0443_),
    .Y(_0469_));
 sky130_fd_sc_hs__clkbuf_8 _4590_ (.A(_0469_),
    .X(_0470_));
 sky130_fd_sc_hs__nor2_2 _4591_ (.A(_0442_),
    .B(_0470_),
    .Y(_2275_));
 sky130_fd_sc_hs__nor2_2 _4592_ (.A(_0460_),
    .B(_0466_),
    .Y(_2274_));
 sky130_fd_sc_hs__mux2i_4 _4593_ (.A0(net180),
    .A1(net166),
    .S(_0439_),
    .Y(_0471_));
 sky130_fd_sc_hs__buf_4 _4594_ (.A(_0471_),
    .X(_0472_));
 sky130_fd_sc_hs__nor2_1 _4595_ (.A(_0445_),
    .B(_0472_),
    .Y(_3731_));
 sky130_fd_sc_hs__mux2i_4 _4596_ (.A0(net135),
    .A1(net149),
    .S(_0443_),
    .Y(_0473_));
 sky130_fd_sc_hs__clkbuf_8 _4597_ (.A(_0473_),
    .X(_0474_));
 sky130_fd_sc_hs__nor2_2 _4598_ (.A(_0442_),
    .B(_0474_),
    .Y(_2292_));
 sky130_fd_sc_hs__nor2_2 _4599_ (.A(_0460_),
    .B(_0470_),
    .Y(_2291_));
 sky130_fd_sc_hs__nor2_1 _4600_ (.A(_0453_),
    .B(_0466_),
    .Y(_2298_));
 sky130_fd_sc_hs__nor2_1 _4601_ (.A(_0456_),
    .B(_0464_),
    .Y(_2297_));
 sky130_fd_sc_hs__nor2_1 _4602_ (.A(_0458_),
    .B(_0468_),
    .Y(_2296_));
 sky130_fd_sc_hs__nor2_1 _4603_ (.A(_0462_),
    .B(_0472_),
    .Y(_3741_));
 sky130_fd_sc_hs__mux2i_4 _4604_ (.A0(net181),
    .A1(net167),
    .S(_0439_),
    .Y(_0475_));
 sky130_fd_sc_hs__clkbuf_8 _4605_ (.A(_0475_),
    .X(_0476_));
 sky130_fd_sc_hs__nor2_1 _4606_ (.A(_0445_),
    .B(_0476_),
    .Y(_3740_));
 sky130_fd_sc_hs__inv_1 _4607_ (.A(_2312_),
    .Y(_2309_));
 sky130_fd_sc_hs__mux2i_4 _4608_ (.A0(net136),
    .A1(net150),
    .S(_0443_),
    .Y(_0477_));
 sky130_fd_sc_hs__clkbuf_8 _4609_ (.A(_0477_),
    .X(_0478_));
 sky130_fd_sc_hs__nor2_2 _4610_ (.A(_0442_),
    .B(_0478_),
    .Y(_2314_));
 sky130_fd_sc_hs__nor2_1 _4611_ (.A(_0460_),
    .B(_0474_),
    .Y(_2313_));
 sky130_fd_sc_hs__nor2_1 _4612_ (.A(_0453_),
    .B(_0470_),
    .Y(_2320_));
 sky130_fd_sc_hs__nor2_1 _4613_ (.A(_0464_),
    .B(_0466_),
    .Y(_2319_));
 sky130_fd_sc_hs__nor2_1 _4614_ (.A(_0456_),
    .B(_0468_),
    .Y(_2318_));
 sky130_fd_sc_hs__nor2_1 _4615_ (.A(_0458_),
    .B(_0472_),
    .Y(_2330_));
 sky130_fd_sc_hs__nor2_1 _4616_ (.A(_0462_),
    .B(_0476_),
    .Y(_2329_));
 sky130_fd_sc_hs__mux2i_4 _4617_ (.A0(net182),
    .A1(net168),
    .S(_0439_),
    .Y(_0479_));
 sky130_fd_sc_hs__buf_4 _4618_ (.A(_0479_),
    .X(_0480_));
 sky130_fd_sc_hs__nor2_2 _4619_ (.A(_0445_),
    .B(_0480_),
    .Y(_2328_));
 sky130_fd_sc_hs__inv_1 _4620_ (.A(_2342_),
    .Y(_2339_));
 sky130_fd_sc_hs__mux2i_4 _4621_ (.A0(net137),
    .A1(net151),
    .S(_0443_),
    .Y(_0481_));
 sky130_fd_sc_hs__clkbuf_8 _4622_ (.A(_0481_),
    .X(_0482_));
 sky130_fd_sc_hs__nor2_2 _4623_ (.A(_0442_),
    .B(_0482_),
    .Y(_2349_));
 sky130_fd_sc_hs__nor2_1 _4624_ (.A(_0460_),
    .B(_0478_),
    .Y(_2348_));
 sky130_fd_sc_hs__nor2_1 _4625_ (.A(_0453_),
    .B(_0474_),
    .Y(_2355_));
 sky130_fd_sc_hs__nor2_1 _4626_ (.A(_0464_),
    .B(_0470_),
    .Y(_2354_));
 sky130_fd_sc_hs__nor2_1 _4627_ (.A(_0466_),
    .B(_0468_),
    .Y(_2353_));
 sky130_fd_sc_hs__nor2_1 _4628_ (.A(_0456_),
    .B(_0472_),
    .Y(_2365_));
 sky130_fd_sc_hs__nor2_1 _4629_ (.A(_0458_),
    .B(_0476_),
    .Y(_2364_));
 sky130_fd_sc_hs__nor2_1 _4630_ (.A(_0462_),
    .B(_0480_),
    .Y(_2363_));
 sky130_fd_sc_hs__mux2i_4 _4631_ (.A0(net183),
    .A1(net169),
    .S(_0439_),
    .Y(_0483_));
 sky130_fd_sc_hs__buf_4 _4632_ (.A(_0483_),
    .X(_0484_));
 sky130_fd_sc_hs__nor2_4 _4633_ (.A(_0445_),
    .B(_0484_),
    .Y(_3757_));
 sky130_fd_sc_hs__mux2i_4 _4634_ (.A0(net138),
    .A1(net152),
    .S(_0454_),
    .Y(_0485_));
 sky130_fd_sc_hs__clkbuf_8 _4635_ (.A(_0485_),
    .X(_0486_));
 sky130_fd_sc_hs__nor2_1 _4636_ (.A(_0442_),
    .B(_0486_),
    .Y(_2377_));
 sky130_fd_sc_hs__nor2_1 _4637_ (.A(_0453_),
    .B(_0478_),
    .Y(_2383_));
 sky130_fd_sc_hs__nor2_1 _4638_ (.A(_0464_),
    .B(_0474_),
    .Y(_2382_));
 sky130_fd_sc_hs__nor2_1 _4639_ (.A(_0468_),
    .B(_0470_),
    .Y(_2381_));
 sky130_fd_sc_hs__nor2_1 _4640_ (.A(_0466_),
    .B(_0472_),
    .Y(_2393_));
 sky130_fd_sc_hs__nor2_1 _4641_ (.A(_0456_),
    .B(_0476_),
    .Y(_2392_));
 sky130_fd_sc_hs__nor2_1 _4642_ (.A(_0458_),
    .B(_0480_),
    .Y(_2391_));
 sky130_fd_sc_hs__nor2_1 _4643_ (.A(_0462_),
    .B(_0484_),
    .Y(_3768_));
 sky130_fd_sc_hs__mux2i_4 _4644_ (.A0(net184),
    .A1(net170),
    .S(_0439_),
    .Y(_0487_));
 sky130_fd_sc_hs__buf_4 _4645_ (.A(_0487_),
    .X(_0488_));
 sky130_fd_sc_hs__nor2_1 _4646_ (.A(_0445_),
    .B(_0488_),
    .Y(_3767_));
 sky130_fd_sc_hs__inv_1 _4647_ (.A(_2407_),
    .Y(_2404_));
 sky130_fd_sc_hs__mux2i_4 _4648_ (.A0(net139),
    .A1(net122),
    .S(_0454_),
    .Y(_0489_));
 sky130_fd_sc_hs__clkbuf_8 _4649_ (.A(_0489_),
    .X(_0490_));
 sky130_fd_sc_hs__nor2_1 _4650_ (.A(_0442_),
    .B(_0490_),
    .Y(_2409_));
 sky130_fd_sc_hs__nor2_1 _4651_ (.A(_0453_),
    .B(_0482_),
    .Y(_2415_));
 sky130_fd_sc_hs__nor2_1 _4652_ (.A(_0464_),
    .B(_0478_),
    .Y(_2414_));
 sky130_fd_sc_hs__nor2_1 _4653_ (.A(_0468_),
    .B(_0474_),
    .Y(_2413_));
 sky130_fd_sc_hs__nor2_1 _4654_ (.A(_0470_),
    .B(_0472_),
    .Y(_2425_));
 sky130_fd_sc_hs__nor2_1 _4655_ (.A(_0466_),
    .B(_0476_),
    .Y(_2424_));
 sky130_fd_sc_hs__nor2_1 _4656_ (.A(_0456_),
    .B(_0480_),
    .Y(_2423_));
 sky130_fd_sc_hs__nor2_1 _4657_ (.A(_0458_),
    .B(_0484_),
    .Y(_2437_));
 sky130_fd_sc_hs__nor2_1 _4658_ (.A(_0462_),
    .B(_0488_),
    .Y(_2436_));
 sky130_fd_sc_hs__mux2i_4 _4659_ (.A0(net154),
    .A1(net171),
    .S(_0440_),
    .Y(_0491_));
 sky130_fd_sc_hs__buf_4 _4660_ (.A(_0491_),
    .X(_0492_));
 sky130_fd_sc_hs__nor2_2 _4661_ (.A(_0444_),
    .B(_0492_),
    .Y(_2435_));
 sky130_fd_sc_hs__mux2i_4 _4662_ (.A0(net140),
    .A1(net123),
    .S(_0454_),
    .Y(_0493_));
 sky130_fd_sc_hs__buf_4 _4663_ (.A(_0493_),
    .X(_0494_));
 sky130_fd_sc_hs__nor2_1 _4664_ (.A(_0442_),
    .B(_0494_),
    .Y(_2447_));
 sky130_fd_sc_hs__nor2_1 _4665_ (.A(_0453_),
    .B(_0486_),
    .Y(_2453_));
 sky130_fd_sc_hs__nor2_1 _4666_ (.A(_0464_),
    .B(_0482_),
    .Y(_2452_));
 sky130_fd_sc_hs__nor2_1 _4667_ (.A(_0468_),
    .B(_0478_),
    .Y(_2451_));
 sky130_fd_sc_hs__nor2_1 _4668_ (.A(_0472_),
    .B(_0474_),
    .Y(_2463_));
 sky130_fd_sc_hs__nor2_1 _4669_ (.A(_0470_),
    .B(_0476_),
    .Y(_2462_));
 sky130_fd_sc_hs__nor2_1 _4670_ (.A(_0466_),
    .B(_0480_),
    .Y(_2461_));
 sky130_fd_sc_hs__nor2_1 _4671_ (.A(_0456_),
    .B(_0484_),
    .Y(_2475_));
 sky130_fd_sc_hs__nor2_1 _4672_ (.A(_0458_),
    .B(_0488_),
    .Y(_2474_));
 sky130_fd_sc_hs__nor2_1 _4673_ (.A(_0462_),
    .B(_0492_),
    .Y(_2473_));
 sky130_fd_sc_hs__mux2i_4 _4674_ (.A0(net155),
    .A1(net172),
    .S(_0440_),
    .Y(_0495_));
 sky130_fd_sc_hs__buf_4 _4675_ (.A(_0495_),
    .X(_0496_));
 sky130_fd_sc_hs__nor2_2 _4676_ (.A(_0444_),
    .B(_0496_),
    .Y(_2478_));
 sky130_fd_sc_hs__mux2i_4 _4677_ (.A0(net141),
    .A1(net124),
    .S(_0454_),
    .Y(_0497_));
 sky130_fd_sc_hs__buf_4 _4678_ (.A(_0497_),
    .X(_0498_));
 sky130_fd_sc_hs__nor2_1 _4679_ (.A(_0441_),
    .B(_0498_),
    .Y(_2492_));
 sky130_fd_sc_hs__nor2_1 _4680_ (.A(_0453_),
    .B(_0490_),
    .Y(_2498_));
 sky130_fd_sc_hs__nor2_1 _4681_ (.A(_0464_),
    .B(_0486_),
    .Y(_2497_));
 sky130_fd_sc_hs__nor2_1 _4682_ (.A(_0468_),
    .B(_0482_),
    .Y(_2496_));
 sky130_fd_sc_hs__nor2_1 _4683_ (.A(_0472_),
    .B(_0478_),
    .Y(_2508_));
 sky130_fd_sc_hs__nor2_1 _4684_ (.A(_0474_),
    .B(_0476_),
    .Y(_2507_));
 sky130_fd_sc_hs__nor2_1 _4685_ (.A(_0470_),
    .B(_0480_),
    .Y(_2506_));
 sky130_fd_sc_hs__nor2_1 _4686_ (.A(_0466_),
    .B(_0484_),
    .Y(_2520_));
 sky130_fd_sc_hs__nor2_1 _4687_ (.A(_0456_),
    .B(_0488_),
    .Y(_2519_));
 sky130_fd_sc_hs__nor2_1 _4688_ (.A(_0458_),
    .B(_0492_),
    .Y(_2518_));
 sky130_fd_sc_hs__nor2_1 _4689_ (.A(_0462_),
    .B(_0496_),
    .Y(_3794_));
 sky130_fd_sc_hs__mux2i_4 _4690_ (.A0(net156),
    .A1(net173),
    .S(_0440_),
    .Y(_0499_));
 sky130_fd_sc_hs__buf_4 _4691_ (.A(_0499_),
    .X(_0500_));
 sky130_fd_sc_hs__nor2_1 _4692_ (.A(_0444_),
    .B(_0500_),
    .Y(_3793_));
 sky130_fd_sc_hs__mux2i_4 _4693_ (.A0(net142),
    .A1(net125),
    .S(_0454_),
    .Y(_0501_));
 sky130_fd_sc_hs__buf_4 _4694_ (.A(_0501_),
    .X(_0502_));
 sky130_fd_sc_hs__nor2_1 _4695_ (.A(_0441_),
    .B(_0502_),
    .Y(_2538_));
 sky130_fd_sc_hs__nor2_1 _4696_ (.A(_0452_),
    .B(_0494_),
    .Y(_2544_));
 sky130_fd_sc_hs__nor2_1 _4697_ (.A(_0464_),
    .B(_0490_),
    .Y(_2543_));
 sky130_fd_sc_hs__nor2_1 _4698_ (.A(_0468_),
    .B(_0486_),
    .Y(_2542_));
 sky130_fd_sc_hs__nor2_1 _4699_ (.A(_0472_),
    .B(_0482_),
    .Y(_2554_));
 sky130_fd_sc_hs__nor2_1 _4700_ (.A(_0476_),
    .B(_0478_),
    .Y(_2553_));
 sky130_fd_sc_hs__nor2_1 _4701_ (.A(_0474_),
    .B(_0480_),
    .Y(_2552_));
 sky130_fd_sc_hs__nor2_1 _4702_ (.A(_0470_),
    .B(_0484_),
    .Y(_2566_));
 sky130_fd_sc_hs__nor2_1 _4703_ (.A(_0466_),
    .B(_0488_),
    .Y(_2565_));
 sky130_fd_sc_hs__nor2_2 _4704_ (.A(_0456_),
    .B(_0492_),
    .Y(_2564_));
 sky130_fd_sc_hs__nor2_1 _4705_ (.A(_0458_),
    .B(_0496_),
    .Y(_2571_));
 sky130_fd_sc_hs__nor2_1 _4706_ (.A(_0462_),
    .B(_0500_),
    .Y(_2570_));
 sky130_fd_sc_hs__mux2i_4 _4707_ (.A0(net157),
    .A1(net174),
    .S(_0440_),
    .Y(_0503_));
 sky130_fd_sc_hs__buf_4 _4708_ (.A(_0503_),
    .X(_0504_));
 sky130_fd_sc_hs__nor2_2 _4709_ (.A(_0444_),
    .B(_0504_),
    .Y(_2569_));
 sky130_fd_sc_hs__mux2i_4 _4710_ (.A0(net144),
    .A1(net126),
    .S(_0454_),
    .Y(_0505_));
 sky130_fd_sc_hs__buf_4 _4711_ (.A(_0505_),
    .X(_0506_));
 sky130_fd_sc_hs__nor2_1 _4712_ (.A(_0441_),
    .B(_0506_),
    .Y(_2593_));
 sky130_fd_sc_hs__nor2_1 _4713_ (.A(_0452_),
    .B(_0498_),
    .Y(_2599_));
 sky130_fd_sc_hs__nor2_1 _4714_ (.A(_0463_),
    .B(_0494_),
    .Y(_2598_));
 sky130_fd_sc_hs__nor2_2 _4715_ (.A(_0468_),
    .B(_0490_),
    .Y(_2597_));
 sky130_fd_sc_hs__nor2_1 _4716_ (.A(_0472_),
    .B(_0486_),
    .Y(_2609_));
 sky130_fd_sc_hs__nor2_1 _4717_ (.A(_0476_),
    .B(_0482_),
    .Y(_2608_));
 sky130_fd_sc_hs__nor2_1 _4718_ (.A(_0478_),
    .B(_0480_),
    .Y(_2607_));
 sky130_fd_sc_hs__nor2_1 _4719_ (.A(_0474_),
    .B(_0484_),
    .Y(_2621_));
 sky130_fd_sc_hs__nor2_1 _4720_ (.A(_0470_),
    .B(_0488_),
    .Y(_2620_));
 sky130_fd_sc_hs__nor2_2 _4721_ (.A(_0465_),
    .B(_0492_),
    .Y(_2619_));
 sky130_fd_sc_hs__nor2_1 _4722_ (.A(_0455_),
    .B(_0496_),
    .Y(_2626_));
 sky130_fd_sc_hs__nor2_2 _4723_ (.A(_0457_),
    .B(_0500_),
    .Y(_2625_));
 sky130_fd_sc_hs__nor2_1 _4724_ (.A(_0461_),
    .B(_0504_),
    .Y(_2624_));
 sky130_fd_sc_hs__mux2i_4 _4725_ (.A0(net158),
    .A1(net176),
    .S(_0440_),
    .Y(_0507_));
 sky130_fd_sc_hs__buf_4 _4726_ (.A(_0507_),
    .X(_0508_));
 sky130_fd_sc_hs__nor2_1 _4727_ (.A(_0444_),
    .B(_0508_),
    .Y(_3807_));
 sky130_fd_sc_hs__inv_1 _4728_ (.A(_2649_),
    .Y(_2645_));
 sky130_fd_sc_hs__mux2i_4 _4729_ (.A0(net145),
    .A1(net127),
    .S(_0454_),
    .Y(_0509_));
 sky130_fd_sc_hs__buf_4 _4730_ (.A(_0509_),
    .X(_0510_));
 sky130_fd_sc_hs__nor2_1 _4731_ (.A(_0441_),
    .B(_0510_),
    .Y(_2651_));
 sky130_fd_sc_hs__nor2_1 _4732_ (.A(_0452_),
    .B(_0502_),
    .Y(_2657_));
 sky130_fd_sc_hs__nor2_1 _4733_ (.A(_0463_),
    .B(_0498_),
    .Y(_2656_));
 sky130_fd_sc_hs__nor2_1 _4734_ (.A(_0467_),
    .B(_0494_),
    .Y(_2655_));
 sky130_fd_sc_hs__nor2_1 _4735_ (.A(_0471_),
    .B(_0490_),
    .Y(_2667_));
 sky130_fd_sc_hs__nor2_1 _4736_ (.A(_0476_),
    .B(_0486_),
    .Y(_2666_));
 sky130_fd_sc_hs__nor2_1 _4737_ (.A(_0480_),
    .B(_0482_),
    .Y(_2665_));
 sky130_fd_sc_hs__nor2_1 _4738_ (.A(_0478_),
    .B(_0484_),
    .Y(_2679_));
 sky130_fd_sc_hs__nor2_1 _4739_ (.A(_0474_),
    .B(_0488_),
    .Y(_2678_));
 sky130_fd_sc_hs__nor2_1 _4740_ (.A(_0469_),
    .B(_0492_),
    .Y(_2677_));
 sky130_fd_sc_hs__nor2_1 _4741_ (.A(_0465_),
    .B(_0496_),
    .Y(_2684_));
 sky130_fd_sc_hs__nor2_1 _4742_ (.A(_0455_),
    .B(_0500_),
    .Y(_2683_));
 sky130_fd_sc_hs__nor2_1 _4743_ (.A(_0457_),
    .B(_0504_),
    .Y(_2682_));
 sky130_fd_sc_hs__nor2_1 _4744_ (.A(_0461_),
    .B(_0508_),
    .Y(_3815_));
 sky130_fd_sc_hs__mux2i_4 _4745_ (.A0(net159),
    .A1(net177),
    .S(_0440_),
    .Y(_0511_));
 sky130_fd_sc_hs__buf_4 _4746_ (.A(_0511_),
    .X(_0512_));
 sky130_fd_sc_hs__nor2_1 _4747_ (.A(_0444_),
    .B(_0512_),
    .Y(_3814_));
 sky130_fd_sc_hs__inv_1 _4748_ (.A(_2702_),
    .Y(_2699_));
 sky130_fd_sc_hs__a22o_4 _4749_ (.A1(_0081_),
    .A2(net114),
    .B1(_0086_),
    .B2(_0436_),
    .X(_2704_));
 sky130_fd_sc_hs__and2_2 _4750_ (.A(net145),
    .B(net188),
    .X(_0513_));
 sky130_fd_sc_hs__nand2b_4 _4751_ (.A_N(_0443_),
    .B(_0513_),
    .Y(_0514_));
 sky130_fd_sc_hs__nor2_8 _4752_ (.A(_0441_),
    .B(_0514_),
    .Y(_2703_));
 sky130_fd_sc_hs__clkinv_8 _4753_ (.A(_2703_),
    .Y(_2779_));
 sky130_fd_sc_hs__nor2_1 _4754_ (.A(_0460_),
    .B(_0510_),
    .Y(_2710_));
 sky130_fd_sc_hs__nor2_1 _4755_ (.A(_0452_),
    .B(_0506_),
    .Y(_2709_));
 sky130_fd_sc_hs__nor2_1 _4756_ (.A(_0463_),
    .B(_0502_),
    .Y(_2708_));
 sky130_fd_sc_hs__nor2_1 _4757_ (.A(_0467_),
    .B(_0498_),
    .Y(_2720_));
 sky130_fd_sc_hs__nor2_1 _4758_ (.A(_0471_),
    .B(_0494_),
    .Y(_2719_));
 sky130_fd_sc_hs__nor2_1 _4759_ (.A(_0475_),
    .B(_0490_),
    .Y(_2718_));
 sky130_fd_sc_hs__nor2_2 _4760_ (.A(_0480_),
    .B(_0486_),
    .Y(_2732_));
 sky130_fd_sc_hs__nor2_1 _4761_ (.A(_0482_),
    .B(_0484_),
    .Y(_2731_));
 sky130_fd_sc_hs__nor2_1 _4762_ (.A(_0478_),
    .B(_0488_),
    .Y(_2730_));
 sky130_fd_sc_hs__nor2_1 _4763_ (.A(_0473_),
    .B(_0492_),
    .Y(_2737_));
 sky130_fd_sc_hs__nor2_1 _4764_ (.A(_0469_),
    .B(_0496_),
    .Y(_2736_));
 sky130_fd_sc_hs__nor2_1 _4765_ (.A(_0465_),
    .B(_0500_),
    .Y(_2735_));
 sky130_fd_sc_hs__nor2_1 _4766_ (.A(_0455_),
    .B(_0504_),
    .Y(_2751_));
 sky130_fd_sc_hs__nor2_1 _4767_ (.A(_0457_),
    .B(_0508_),
    .Y(_2750_));
 sky130_fd_sc_hs__nor2_2 _4768_ (.A(_0461_),
    .B(_0512_),
    .Y(_2749_));
 sky130_fd_sc_hs__inv_1 _4769_ (.A(_2773_),
    .Y(_2770_));
 sky130_fd_sc_hs__nand2_2 _4770_ (.A(_0081_),
    .B(net115),
    .Y(_0515_));
 sky130_fd_sc_hs__nand2_1 _4771_ (.A(_0446_),
    .B(_0086_),
    .Y(_0516_));
 sky130_fd_sc_hs__nand2_4 _4772_ (.A(_0515_),
    .B(_0516_),
    .Y(_2775_));
 sky130_fd_sc_hs__nor2_8 _4773_ (.A(_0459_),
    .B(_0514_),
    .Y(_2774_));
 sky130_fd_sc_hs__nor2_1 _4774_ (.A(_0452_),
    .B(_0510_),
    .Y(_2782_));
 sky130_fd_sc_hs__nor2_1 _4775_ (.A(_0463_),
    .B(_0506_),
    .Y(_2781_));
 sky130_fd_sc_hs__nor2_1 _4776_ (.A(_0467_),
    .B(_0502_),
    .Y(_2780_));
 sky130_fd_sc_hs__nor2_1 _4777_ (.A(_0471_),
    .B(_0498_),
    .Y(_2792_));
 sky130_fd_sc_hs__nor2_1 _4778_ (.A(_0475_),
    .B(_0494_),
    .Y(_2791_));
 sky130_fd_sc_hs__nor2_1 _4779_ (.A(_0479_),
    .B(_0490_),
    .Y(_2790_));
 sky130_fd_sc_hs__nor2_1 _4780_ (.A(_0484_),
    .B(_0486_),
    .Y(_2804_));
 sky130_fd_sc_hs__nor2_2 _4781_ (.A(_0482_),
    .B(_0488_),
    .Y(_2803_));
 sky130_fd_sc_hs__nor2_1 _4782_ (.A(_0477_),
    .B(_0492_),
    .Y(_2802_));
 sky130_fd_sc_hs__nor2_1 _4783_ (.A(_0473_),
    .B(_0496_),
    .Y(_2809_));
 sky130_fd_sc_hs__nor2_1 _4784_ (.A(_0469_),
    .B(_0500_),
    .Y(_2808_));
 sky130_fd_sc_hs__nor2_1 _4785_ (.A(_0465_),
    .B(_0504_),
    .Y(_2807_));
 sky130_fd_sc_hs__nor2_1 _4786_ (.A(_0455_),
    .B(_0508_),
    .Y(_2823_));
 sky130_fd_sc_hs__nor2_1 _4787_ (.A(_0457_),
    .B(_0512_),
    .Y(_2822_));
 sky130_fd_sc_hs__and2_1 _4788_ (.A(net177),
    .B(net189),
    .X(_0517_));
 sky130_fd_sc_hs__and2_4 _4789_ (.A(_0440_),
    .B(_0517_),
    .X(_0518_));
 sky130_fd_sc_hs__clkbuf_8 _4790_ (.A(_0518_),
    .X(_2705_));
 sky130_fd_sc_hs__and2_1 _4791_ (.A(_0461_),
    .B(_2705_),
    .X(_2821_));
 sky130_fd_sc_hs__buf_8 _4792_ (.A(_0514_),
    .X(_0519_));
 sky130_fd_sc_hs__nor2_4 _4793_ (.A(_0452_),
    .B(_0519_),
    .Y(_2844_));
 sky130_fd_sc_hs__nor2_1 _4794_ (.A(_0463_),
    .B(_0510_),
    .Y(_2843_));
 sky130_fd_sc_hs__nor2_1 _4795_ (.A(_0467_),
    .B(_0506_),
    .Y(_2842_));
 sky130_fd_sc_hs__nor2_1 _4796_ (.A(_0471_),
    .B(_0502_),
    .Y(_2854_));
 sky130_fd_sc_hs__nor2_1 _4797_ (.A(_0475_),
    .B(_0498_),
    .Y(_2853_));
 sky130_fd_sc_hs__nor2_1 _4798_ (.A(_0479_),
    .B(_0494_),
    .Y(_2852_));
 sky130_fd_sc_hs__nor2_2 _4799_ (.A(_0483_),
    .B(_0490_),
    .Y(_2866_));
 sky130_fd_sc_hs__nor2_2 _4800_ (.A(_0486_),
    .B(_0488_),
    .Y(_2865_));
 sky130_fd_sc_hs__nor2_1 _4801_ (.A(_0481_),
    .B(_0492_),
    .Y(_2864_));
 sky130_fd_sc_hs__nor2_1 _4802_ (.A(_0477_),
    .B(_0496_),
    .Y(_2871_));
 sky130_fd_sc_hs__nor2_1 _4803_ (.A(_0473_),
    .B(_0500_),
    .Y(_2870_));
 sky130_fd_sc_hs__nor2_1 _4804_ (.A(_0469_),
    .B(_0504_),
    .Y(_2869_));
 sky130_fd_sc_hs__nor2_1 _4805_ (.A(_0465_),
    .B(_0508_),
    .Y(_2885_));
 sky130_fd_sc_hs__nor2_1 _4806_ (.A(_0455_),
    .B(_0512_),
    .Y(_2884_));
 sky130_fd_sc_hs__and2_1 _4807_ (.A(_0457_),
    .B(_2705_),
    .X(_2883_));
 sky130_fd_sc_hs__nor2_4 _4808_ (.A(_0463_),
    .B(_0519_),
    .Y(_2907_));
 sky130_fd_sc_hs__nor2_1 _4809_ (.A(_0467_),
    .B(_0510_),
    .Y(_2906_));
 sky130_fd_sc_hs__nor2_1 _4810_ (.A(_0471_),
    .B(_0506_),
    .Y(_2917_));
 sky130_fd_sc_hs__nor2_1 _4811_ (.A(_0475_),
    .B(_0502_),
    .Y(_2916_));
 sky130_fd_sc_hs__nor2_1 _4812_ (.A(_0479_),
    .B(_0498_),
    .Y(_2915_));
 sky130_fd_sc_hs__nor2_1 _4813_ (.A(_0483_),
    .B(_0494_),
    .Y(_2929_));
 sky130_fd_sc_hs__nor2_2 _4814_ (.A(_0487_),
    .B(_0490_),
    .Y(_2928_));
 sky130_fd_sc_hs__nor2_2 _4815_ (.A(_0485_),
    .B(_0492_),
    .Y(_2927_));
 sky130_fd_sc_hs__nor2_1 _4816_ (.A(_0481_),
    .B(_0496_),
    .Y(_2934_));
 sky130_fd_sc_hs__nor2_1 _4817_ (.A(_0477_),
    .B(_0500_),
    .Y(_2933_));
 sky130_fd_sc_hs__nor2_1 _4818_ (.A(_0473_),
    .B(_0504_),
    .Y(_2932_));
 sky130_fd_sc_hs__nor2_1 _4819_ (.A(_0469_),
    .B(_0508_),
    .Y(_2948_));
 sky130_fd_sc_hs__nor2_1 _4820_ (.A(_0465_),
    .B(_0512_),
    .Y(_2947_));
 sky130_fd_sc_hs__and2_1 _4821_ (.A(_0455_),
    .B(_2705_),
    .X(_2946_));
 sky130_fd_sc_hs__nor2_1 _4822_ (.A(_0467_),
    .B(_0519_),
    .Y(_2970_));
 sky130_fd_sc_hs__nor2_1 _4823_ (.A(_0471_),
    .B(_0510_),
    .Y(_2980_));
 sky130_fd_sc_hs__nor2_1 _4824_ (.A(_0475_),
    .B(_0506_),
    .Y(_2979_));
 sky130_fd_sc_hs__nor2_1 _4825_ (.A(_0479_),
    .B(_0502_),
    .Y(_2978_));
 sky130_fd_sc_hs__nor2_1 _4826_ (.A(_0483_),
    .B(_0498_),
    .Y(_2992_));
 sky130_fd_sc_hs__nor2_1 _4827_ (.A(_0487_),
    .B(_0494_),
    .Y(_2991_));
 sky130_fd_sc_hs__nor2_1 _4828_ (.A(_0489_),
    .B(_0491_),
    .Y(_2990_));
 sky130_fd_sc_hs__nor2_1 _4829_ (.A(_0485_),
    .B(_0496_),
    .Y(_2997_));
 sky130_fd_sc_hs__nor2_1 _4830_ (.A(_0481_),
    .B(_0500_),
    .Y(_2996_));
 sky130_fd_sc_hs__nor2_1 _4831_ (.A(_0477_),
    .B(_0504_),
    .Y(_2995_));
 sky130_fd_sc_hs__nor2_1 _4832_ (.A(_0473_),
    .B(_0508_),
    .Y(_3011_));
 sky130_fd_sc_hs__nor2_1 _4833_ (.A(_0469_),
    .B(_0512_),
    .Y(_3010_));
 sky130_fd_sc_hs__and2_1 _4834_ (.A(_0465_),
    .B(_2705_),
    .X(_3009_));
 sky130_fd_sc_hs__nor2_4 _4835_ (.A(_0471_),
    .B(_0519_),
    .Y(_3039_));
 sky130_fd_sc_hs__nor2_1 _4836_ (.A(_0475_),
    .B(_0510_),
    .Y(_3038_));
 sky130_fd_sc_hs__nor2_1 _4837_ (.A(_0479_),
    .B(_0506_),
    .Y(_3037_));
 sky130_fd_sc_hs__nor2_1 _4838_ (.A(_0483_),
    .B(_0502_),
    .Y(_3051_));
 sky130_fd_sc_hs__nor2_1 _4839_ (.A(_0487_),
    .B(_0498_),
    .Y(_3050_));
 sky130_fd_sc_hs__nor2_2 _4840_ (.A(_0491_),
    .B(_0494_),
    .Y(_3049_));
 sky130_fd_sc_hs__nor2_1 _4841_ (.A(_0489_),
    .B(_0495_),
    .Y(_3056_));
 sky130_fd_sc_hs__nor2_2 _4842_ (.A(_0485_),
    .B(_0500_),
    .Y(_3055_));
 sky130_fd_sc_hs__nor2_1 _4843_ (.A(_0481_),
    .B(_0504_),
    .Y(_3054_));
 sky130_fd_sc_hs__nor2_1 _4844_ (.A(_0477_),
    .B(_0508_),
    .Y(_3070_));
 sky130_fd_sc_hs__nor2_1 _4845_ (.A(_0473_),
    .B(_0512_),
    .Y(_3069_));
 sky130_fd_sc_hs__and2_1 _4846_ (.A(_0469_),
    .B(_2705_),
    .X(_3068_));
 sky130_fd_sc_hs__clkbuf_16 _4847_ (.A(imd_val_q_i[56]),
    .X(_0520_));
 sky130_fd_sc_hs__clkbuf_8 _4848_ (.A(_0085_),
    .X(_0521_));
 sky130_fd_sc_hs__inv_1 _4849_ (.A(net188),
    .Y(_0522_));
 sky130_fd_sc_hs__inv_2 _4850_ (.A(net189),
    .Y(_0523_));
 sky130_fd_sc_hs__a21oi_2 _4851_ (.A1(_0522_),
    .A2(_0523_),
    .B1(_0515_),
    .Y(_0524_));
 sky130_fd_sc_hs__buf_8 _4852_ (.A(_0524_),
    .X(_0525_));
 sky130_fd_sc_hs__a21oi_2 _4853_ (.A1(_0520_),
    .A2(_0521_),
    .B1(_0525_),
    .Y(_3089_));
 sky130_fd_sc_hs__nor2_4 _4854_ (.A(_0475_),
    .B(_0519_),
    .Y(_3096_));
 sky130_fd_sc_hs__nor2_1 _4855_ (.A(_0479_),
    .B(_0510_),
    .Y(_3095_));
 sky130_fd_sc_hs__nor2_1 _4856_ (.A(_0483_),
    .B(_0506_),
    .Y(_3108_));
 sky130_fd_sc_hs__nor2_1 _4857_ (.A(_0487_),
    .B(_0502_),
    .Y(_3107_));
 sky130_fd_sc_hs__nor2_2 _4858_ (.A(_0491_),
    .B(_0498_),
    .Y(_3106_));
 sky130_fd_sc_hs__nor2_1 _4859_ (.A(_0493_),
    .B(_0495_),
    .Y(_3113_));
 sky130_fd_sc_hs__nor2_1 _4860_ (.A(_0489_),
    .B(_0499_),
    .Y(_3112_));
 sky130_fd_sc_hs__nor2_2 _4861_ (.A(_0485_),
    .B(_0504_),
    .Y(_3111_));
 sky130_fd_sc_hs__nor2_1 _4862_ (.A(_0481_),
    .B(_0508_),
    .Y(_3127_));
 sky130_fd_sc_hs__nor2_1 _4863_ (.A(_0477_),
    .B(_0512_),
    .Y(_3126_));
 sky130_fd_sc_hs__and2_1 _4864_ (.A(_0473_),
    .B(_2705_),
    .X(_3125_));
 sky130_fd_sc_hs__buf_8 _4865_ (.A(imd_val_q_i[57]),
    .X(_0526_));
 sky130_fd_sc_hs__a21oi_4 _4866_ (.A1(_0526_),
    .A2(_0521_),
    .B1(_0525_),
    .Y(_3146_));
 sky130_fd_sc_hs__nor2_2 _4867_ (.A(_0479_),
    .B(_0519_),
    .Y(_3153_));
 sky130_fd_sc_hs__nor2_1 _4868_ (.A(_0483_),
    .B(_0510_),
    .Y(_3166_));
 sky130_fd_sc_hs__nor2_1 _4869_ (.A(_0487_),
    .B(_0506_),
    .Y(_3165_));
 sky130_fd_sc_hs__nor2_2 _4870_ (.A(_0491_),
    .B(_0502_),
    .Y(_3164_));
 sky130_fd_sc_hs__nor2_1 _4871_ (.A(_0495_),
    .B(_0497_),
    .Y(_3171_));
 sky130_fd_sc_hs__nor2_1 _4872_ (.A(_0493_),
    .B(_0499_),
    .Y(_3170_));
 sky130_fd_sc_hs__nor2_1 _4873_ (.A(_0489_),
    .B(_0503_),
    .Y(_3169_));
 sky130_fd_sc_hs__nor2_1 _4874_ (.A(_0485_),
    .B(_0508_),
    .Y(_3185_));
 sky130_fd_sc_hs__nor2_1 _4875_ (.A(_0481_),
    .B(_0512_),
    .Y(_3184_));
 sky130_fd_sc_hs__and2_1 _4876_ (.A(_0477_),
    .B(_2705_),
    .X(_3183_));
 sky130_fd_sc_hs__clkbuf_16 _4877_ (.A(imd_val_q_i[58]),
    .X(_0527_));
 sky130_fd_sc_hs__a21oi_4 _4878_ (.A1(_0527_),
    .A2(_0521_),
    .B1(_0525_),
    .Y(_3204_));
 sky130_fd_sc_hs__nor2_4 _4879_ (.A(_0483_),
    .B(_0519_),
    .Y(_3220_));
 sky130_fd_sc_hs__nor2_1 _4880_ (.A(_0487_),
    .B(_0510_),
    .Y(_3219_));
 sky130_fd_sc_hs__nor2_1 _4881_ (.A(_0491_),
    .B(_0506_),
    .Y(_3218_));
 sky130_fd_sc_hs__nor2_1 _4882_ (.A(_0495_),
    .B(_0501_),
    .Y(_3225_));
 sky130_fd_sc_hs__nor2_1 _4883_ (.A(_0497_),
    .B(_0499_),
    .Y(_3224_));
 sky130_fd_sc_hs__nor2_1 _4884_ (.A(_0493_),
    .B(_0503_),
    .Y(_3223_));
 sky130_fd_sc_hs__nor2_1 _4885_ (.A(_0489_),
    .B(_0507_),
    .Y(_3239_));
 sky130_fd_sc_hs__nor2_2 _4886_ (.A(_0485_),
    .B(_0512_),
    .Y(_3238_));
 sky130_fd_sc_hs__and2_1 _4887_ (.A(_0481_),
    .B(_2705_),
    .X(_3237_));
 sky130_fd_sc_hs__o211ai_4 _4888_ (.A1(net188),
    .A2(net189),
    .B1(net115),
    .C1(_0081_),
    .Y(_0528_));
 sky130_fd_sc_hs__buf_8 _4889_ (.A(imd_val_q_i[59]),
    .X(_0529_));
 sky130_fd_sc_hs__nand2_1 _4890_ (.A(_0529_),
    .B(_0086_),
    .Y(_0530_));
 sky130_fd_sc_hs__nand2_2 _4891_ (.A(_0528_),
    .B(_0530_),
    .Y(_3258_));
 sky130_fd_sc_hs__nor2_4 _4892_ (.A(_0487_),
    .B(_0519_),
    .Y(_3269_));
 sky130_fd_sc_hs__nor2_1 _4893_ (.A(_0491_),
    .B(_0509_),
    .Y(_3268_));
 sky130_fd_sc_hs__nor2_1 _4894_ (.A(_0495_),
    .B(_0505_),
    .Y(_3274_));
 sky130_fd_sc_hs__nor2_1 _4895_ (.A(_0499_),
    .B(_0501_),
    .Y(_3273_));
 sky130_fd_sc_hs__nor2_1 _4896_ (.A(_0497_),
    .B(_0503_),
    .Y(_3272_));
 sky130_fd_sc_hs__nor2_1 _4897_ (.A(_0493_),
    .B(_0507_),
    .Y(_3289_));
 sky130_fd_sc_hs__nor2_1 _4898_ (.A(_0489_),
    .B(_0511_),
    .Y(_3288_));
 sky130_fd_sc_hs__and2_1 _4899_ (.A(_0485_),
    .B(_0518_),
    .X(_3287_));
 sky130_fd_sc_hs__nor2_2 _4900_ (.A(_0491_),
    .B(_0519_),
    .Y(_3317_));
 sky130_fd_sc_hs__nor2_1 _4901_ (.A(_0495_),
    .B(_0509_),
    .Y(_3322_));
 sky130_fd_sc_hs__nor2_1 _4902_ (.A(_0499_),
    .B(_0505_),
    .Y(_3321_));
 sky130_fd_sc_hs__nor2_1 _4903_ (.A(_0501_),
    .B(_0503_),
    .Y(_3320_));
 sky130_fd_sc_hs__nor2_1 _4904_ (.A(_0497_),
    .B(_0507_),
    .Y(_3338_));
 sky130_fd_sc_hs__nor2_1 _4905_ (.A(_0493_),
    .B(_0511_),
    .Y(_3337_));
 sky130_fd_sc_hs__and2_1 _4906_ (.A(_0489_),
    .B(_0518_),
    .X(_3336_));
 sky130_fd_sc_hs__nor2_4 _4907_ (.A(_0495_),
    .B(_0519_),
    .Y(_3367_));
 sky130_fd_sc_hs__nor2_1 _4908_ (.A(_0499_),
    .B(_0509_),
    .Y(_3366_));
 sky130_fd_sc_hs__nor2_1 _4909_ (.A(_0503_),
    .B(_0505_),
    .Y(_3365_));
 sky130_fd_sc_hs__nor2_1 _4910_ (.A(_0501_),
    .B(_0507_),
    .Y(_3381_));
 sky130_fd_sc_hs__nor2_1 _4911_ (.A(_0497_),
    .B(_0511_),
    .Y(_3380_));
 sky130_fd_sc_hs__and2_1 _4912_ (.A(_0493_),
    .B(_0518_),
    .X(_3379_));
 sky130_fd_sc_hs__nor2_4 _4913_ (.A(_0499_),
    .B(_0514_),
    .Y(_3408_));
 sky130_fd_sc_hs__nor2_1 _4914_ (.A(_0503_),
    .B(_0509_),
    .Y(_3407_));
 sky130_fd_sc_hs__nor2_1 _4915_ (.A(_0505_),
    .B(_0507_),
    .Y(_3420_));
 sky130_fd_sc_hs__nor2_1 _4916_ (.A(_0501_),
    .B(_0511_),
    .Y(_3419_));
 sky130_fd_sc_hs__and2_1 _4917_ (.A(_0497_),
    .B(_0518_),
    .X(_3418_));
 sky130_fd_sc_hs__nor2_2 _4918_ (.A(_0503_),
    .B(_0514_),
    .Y(_3446_));
 sky130_fd_sc_hs__nor2_1 _4919_ (.A(_0507_),
    .B(_0509_),
    .Y(_3458_));
 sky130_fd_sc_hs__nor2_1 _4920_ (.A(_0505_),
    .B(_0511_),
    .Y(_3457_));
 sky130_fd_sc_hs__and2_1 _4921_ (.A(_0501_),
    .B(_0518_),
    .X(_3456_));
 sky130_fd_sc_hs__nor2_4 _4922_ (.A(_0507_),
    .B(_0514_),
    .Y(_3493_));
 sky130_fd_sc_hs__nor2_1 _4923_ (.A(_0509_),
    .B(_0511_),
    .Y(_3492_));
 sky130_fd_sc_hs__and2_1 _4924_ (.A(_0505_),
    .B(_0518_),
    .X(_3491_));
 sky130_fd_sc_hs__nor2_4 _4925_ (.A(_0511_),
    .B(_0514_),
    .Y(_3523_));
 sky130_fd_sc_hs__and2_1 _4926_ (.A(_0509_),
    .B(_0518_),
    .X(_3522_));
 sky130_fd_sc_hs__and2_1 _4927_ (.A(_0514_),
    .B(_0518_),
    .X(_3551_));
 sky130_fd_sc_hs__clkinv_8 _4928_ (.A(_2774_),
    .Y(_2778_));
 sky130_fd_sc_hs__inv_8 _4929_ (.A(_2972_),
    .Y(_2973_));
 sky130_fd_sc_hs__inv_1 _4930_ (.A(_3485_),
    .Y(_3486_));
 sky130_fd_sc_hs__nor3_4 _4931_ (.A(net214),
    .B(_0264_),
    .C(_0425_),
    .Y(_0531_));
 sky130_fd_sc_hs__buf_4 _4932_ (.A(_0110_),
    .X(_0532_));
 sky130_fd_sc_hs__nand2_1 _4933_ (.A(_0118_),
    .B(_0117_),
    .Y(_0533_));
 sky130_fd_sc_hs__nor2_1 _4934_ (.A(_3570_),
    .B(_0112_),
    .Y(_0534_));
 sky130_fd_sc_hs__nor2b_1 _4935_ (.A(net76),
    .B_N(net77),
    .Y(_0535_));
 sky130_fd_sc_hs__nand2b_1 _4936_ (.A_N(_0534_),
    .B(_0535_),
    .Y(_0536_));
 sky130_fd_sc_hs__buf_4 _4937_ (.A(_0114_),
    .X(_0537_));
 sky130_fd_sc_hs__a21oi_1 _4938_ (.A1(_0533_),
    .A2(_0536_),
    .B1(_0537_),
    .Y(_0538_));
 sky130_fd_sc_hs__nand2b_4 _4939_ (.A_N(net77),
    .B(net76),
    .Y(_0539_));
 sky130_fd_sc_hs__nor2_1 _4940_ (.A(_0537_),
    .B(_3574_),
    .Y(_0540_));
 sky130_fd_sc_hs__a2111oi_1 _4941_ (.A1(_0537_),
    .A2(_0534_),
    .B1(_0539_),
    .C1(_0532_),
    .D1(_0540_),
    .Y(_0541_));
 sky130_fd_sc_hs__a21o_4 _4942_ (.A1(_0532_),
    .A2(_0538_),
    .B1(_0541_),
    .X(_0542_));
 sky130_fd_sc_hs__nand2b_1 _4943_ (.A_N(_0118_),
    .B(_0537_),
    .Y(_0543_));
 sky130_fd_sc_hs__o311ai_2 _4944_ (.A1(_0537_),
    .A2(_3570_),
    .A3(_0112_),
    .B1(_0543_),
    .C1(_0532_),
    .Y(_0544_));
 sky130_fd_sc_hs__nor2b_4 _4945_ (.A(_0110_),
    .B_N(_0114_),
    .Y(_0545_));
 sky130_fd_sc_hs__nand2_1 _4946_ (.A(_3574_),
    .B(_0545_),
    .Y(_0546_));
 sky130_fd_sc_hs__a21oi_4 _4947_ (.A1(_0544_),
    .A2(_0546_),
    .B1(_0539_),
    .Y(_0547_));
 sky130_fd_sc_hs__nor2b_4 _4948_ (.A(_0533_),
    .B_N(_0545_),
    .Y(_0548_));
 sky130_fd_sc_hs__nor3_4 _4949_ (.A(_0542_),
    .B(_0547_),
    .C(_0548_),
    .Y(_0549_));
 sky130_fd_sc_hs__o31a_1 _4950_ (.A1(net214),
    .A2(_0264_),
    .A3(_0425_),
    .B1(_0548_),
    .X(_0550_));
 sky130_fd_sc_hs__nor2_1 _4951_ (.A(_0117_),
    .B(_0535_),
    .Y(_0551_));
 sky130_fd_sc_hs__nand2b_1 _4952_ (.A_N(_0114_),
    .B(_0110_),
    .Y(_0552_));
 sky130_fd_sc_hs__o2bb2ai_2 _4953_ (.A1_N(_0117_),
    .A2_N(_0545_),
    .B1(_0551_),
    .B2(_0552_),
    .Y(_0553_));
 sky130_fd_sc_hs__nand2b_4 _4954_ (.A_N(_0110_),
    .B(_3574_),
    .Y(_0554_));
 sky130_fd_sc_hs__nor2_1 _4955_ (.A(_0539_),
    .B(_0554_),
    .Y(_0555_));
 sky130_fd_sc_hs__a21oi_4 _4956_ (.A1(_0112_),
    .A2(_0553_),
    .B1(_0555_),
    .Y(_0556_));
 sky130_fd_sc_hs__xnor2_4 _4957_ (.A(net34),
    .B(_0556_),
    .Y(_0557_));
 sky130_fd_sc_hs__nand2_2 _4958_ (.A(_3930_),
    .B(_0557_),
    .Y(_0558_));
 sky130_fd_sc_hs__o41a_1 _4959_ (.A1(_3930_),
    .A2(_0404_),
    .A3(_0408_),
    .A4(_0409_),
    .B1(_0558_),
    .X(_0559_));
 sky130_fd_sc_hs__mux2_1 _4960_ (.A0(_0547_),
    .A1(_0542_),
    .S(_0559_),
    .X(_0560_));
 sky130_fd_sc_hs__a211o_4 _4961_ (.A1(_0531_),
    .A2(_0549_),
    .B1(_0550_),
    .C1(_0560_),
    .X(net223));
 sky130_fd_sc_hs__inv_2 _4962_ (.A(net53),
    .Y(_3934_));
 sky130_fd_sc_hs__clkinv_4 _4963_ (.A(net64),
    .Y(_3948_));
 sky130_fd_sc_hs__buf_2 _4964_ (.A(net42),
    .X(_0561_));
 sky130_fd_sc_hs__inv_2 _4965_ (.A(_0561_),
    .Y(_0562_));
 sky130_fd_sc_hs__buf_16 _4966_ (.A(_0562_),
    .X(_0563_));
 sky130_fd_sc_hs__buf_16 _4967_ (.A(_0563_),
    .X(_3933_));
 sky130_fd_sc_hs__clkinv_2 _4968_ (.A(net67),
    .Y(_3954_));
 sky130_fd_sc_hs__inv_2 _4969_ (.A(net68),
    .Y(_3960_));
 sky130_fd_sc_hs__clkinv_8 _4970_ (.A(_0314_),
    .Y(net213));
 sky130_fd_sc_hs__inv_4 _4971_ (.A(_0317_),
    .Y(net218));
 sky130_fd_sc_hs__inv_16 _4972_ (.A(_0374_),
    .Y(net195));
 sky130_fd_sc_hs__nand3_4 _4973_ (.A(_0365_),
    .B(_0366_),
    .C(_0369_),
    .Y(net198));
 sky130_fd_sc_hs__o21bai_2 _4974_ (.A1(_0203_),
    .A2(_0204_),
    .B1_N(_0207_),
    .Y(_0564_));
 sky130_fd_sc_hs__xnor2_4 _4975_ (.A(_0169_),
    .B(_0564_),
    .Y(net200));
 sky130_fd_sc_hs__or2_1 _4976_ (.A(_0444_),
    .B(_0459_),
    .X(_2230_));
 sky130_fd_sc_hs__or2_1 _4977_ (.A(_0459_),
    .B(_0461_),
    .X(_2235_));
 sky130_fd_sc_hs__or2_1 _4978_ (.A(_0461_),
    .B(_0467_),
    .X(_2279_));
 sky130_fd_sc_hs__inv_1 _4979_ (.A(_3771_),
    .Y(_2443_));
 sky130_fd_sc_hs__inv_1 _4980_ (.A(_3779_),
    .Y(_2488_));
 sky130_fd_sc_hs__nand2_1 _4981_ (.A(_0445_),
    .B(_2705_),
    .Y(_2757_));
 sky130_fd_sc_hs__buf_8 _4982_ (.A(imd_val_q_i[60]),
    .X(_0565_));
 sky130_fd_sc_hs__a21oi_4 _4983_ (.A1(_0565_),
    .A2(_0521_),
    .B1(_0525_),
    .Y(_3308_));
 sky130_fd_sc_hs__clkbuf_16 _4984_ (.A(imd_val_q_i[61]),
    .X(_0566_));
 sky130_fd_sc_hs__a21oi_2 _4985_ (.A1(_0566_),
    .A2(_0521_),
    .B1(_0525_),
    .Y(_3357_));
 sky130_fd_sc_hs__a21oi_2 _4986_ (.A1(net111),
    .A2(_0521_),
    .B1(_0525_),
    .Y(_3400_));
 sky130_fd_sc_hs__a21oi_2 _4987_ (.A1(net112),
    .A2(_0521_),
    .B1(_0525_),
    .Y(_3439_));
 sky130_fd_sc_hs__buf_8 _4988_ (.A(imd_val_q_i[64]),
    .X(_0567_));
 sky130_fd_sc_hs__a21oi_4 _4989_ (.A1(_0567_),
    .A2(_0521_),
    .B1(_0525_),
    .Y(_3477_));
 sky130_fd_sc_hs__a21oi_4 _4990_ (.A1(_0382_),
    .A2(_0521_),
    .B1(_0525_),
    .Y(_3513_));
 sky130_fd_sc_hs__a21oi_4 _4991_ (.A1(net114),
    .A2(_0521_),
    .B1(_0525_),
    .Y(_3542_));
 sky130_fd_sc_hs__or2_1 _4992_ (.A(_0441_),
    .B(_0461_),
    .X(_2231_));
 sky130_fd_sc_hs__or2_1 _4993_ (.A(_0441_),
    .B(_0457_),
    .X(_2236_));
 sky130_fd_sc_hs__or2_1 _4994_ (.A(_0457_),
    .B(_0463_),
    .X(_2280_));
 sky130_fd_sc_hs__inv_1 _4995_ (.A(_3817_),
    .Y(_2758_));
 sky130_fd_sc_hs__inv_1 _4996_ (.A(_3260_),
    .Y(_3261_));
 sky130_fd_sc_hs__or2_1 _4997_ (.A(_0452_),
    .B(_0455_),
    .X(_2281_));
 sky130_fd_sc_hs__inv_1 _4998_ (.A(_3374_),
    .Y(_3430_));
 sky130_fd_sc_hs__inv_1 _4999_ (.A(_2369_),
    .Y(_2370_));
 sky130_fd_sc_hs__inv_1 _5000_ (.A(_2397_),
    .Y(_2398_));
 sky130_fd_sc_hs__inv_1 _5001_ (.A(_2445_),
    .Y(_3782_));
 sky130_fd_sc_hs__inv_1 _5002_ (.A(_2490_),
    .Y(_3788_));
 sky130_fd_sc_hs__inv_1 _5003_ (.A(_2583_),
    .Y(_2584_));
 sky130_fd_sc_hs__inv_1 _5004_ (.A(_2638_),
    .Y(_2639_));
 sky130_fd_sc_hs__inv_2 _5005_ (.A(_3091_),
    .Y(_3092_));
 sky130_fd_sc_hs__inv_1 _5006_ (.A(_3148_),
    .Y(_3150_));
 sky130_fd_sc_hs__inv_1 _5007_ (.A(_3206_),
    .Y(_3208_));
 sky130_fd_sc_hs__inv_1 _5008_ (.A(_3263_),
    .Y(_3264_));
 sky130_fd_sc_hs__inv_1 _5009_ (.A(_2249_),
    .Y(_2251_));
 sky130_fd_sc_hs__inv_1 _5010_ (.A(_2258_),
    .Y(_2266_));
 sky130_fd_sc_hs__inv_1 _5011_ (.A(_2263_),
    .Y(_2264_));
 sky130_fd_sc_hs__inv_1 _5012_ (.A(_2278_),
    .Y(_2285_));
 sky130_fd_sc_hs__inv_1 _5013_ (.A(_2295_),
    .Y(_2303_));
 sky130_fd_sc_hs__inv_1 _5014_ (.A(_2300_),
    .Y(_2301_));
 sky130_fd_sc_hs__inv_1 _5015_ (.A(_2317_),
    .Y(_2325_));
 sky130_fd_sc_hs__inv_1 _5016_ (.A(_2322_),
    .Y(_2323_));
 sky130_fd_sc_hs__inv_1 _5017_ (.A(_2335_),
    .Y(_2336_));
 sky130_fd_sc_hs__inv_1 _5018_ (.A(_2352_),
    .Y(_2360_));
 sky130_fd_sc_hs__inv_1 _5019_ (.A(_2357_),
    .Y(_2358_));
 sky130_fd_sc_hs__inv_1 _5020_ (.A(_2380_),
    .Y(_2388_));
 sky130_fd_sc_hs__inv_1 _5021_ (.A(_2385_),
    .Y(_2386_));
 sky130_fd_sc_hs__inv_1 _5022_ (.A(_2412_),
    .Y(_2420_));
 sky130_fd_sc_hs__inv_1 _5023_ (.A(_2417_),
    .Y(_2418_));
 sky130_fd_sc_hs__inv_1 _5024_ (.A(_2427_),
    .Y(_2429_));
 sky130_fd_sc_hs__inv_1 _5025_ (.A(_2450_),
    .Y(_2458_));
 sky130_fd_sc_hs__inv_1 _5026_ (.A(_2455_),
    .Y(_2456_));
 sky130_fd_sc_hs__inv_1 _5027_ (.A(_2465_),
    .Y(_2467_));
 sky130_fd_sc_hs__inv_1 _5028_ (.A(_2484_),
    .Y(_2485_));
 sky130_fd_sc_hs__inv_1 _5029_ (.A(_2495_),
    .Y(_2503_));
 sky130_fd_sc_hs__inv_1 _5030_ (.A(_2500_),
    .Y(_2501_));
 sky130_fd_sc_hs__inv_1 _5031_ (.A(_2510_),
    .Y(_2512_));
 sky130_fd_sc_hs__inv_1 _5032_ (.A(_2522_),
    .Y(_2525_));
 sky130_fd_sc_hs__inv_1 _5033_ (.A(_2541_),
    .Y(_2549_));
 sky130_fd_sc_hs__inv_1 _5034_ (.A(_2546_),
    .Y(_2547_));
 sky130_fd_sc_hs__inv_1 _5035_ (.A(_2556_),
    .Y(_2558_));
 sky130_fd_sc_hs__inv_1 _5036_ (.A(_2568_),
    .Y(_2576_));
 sky130_fd_sc_hs__inv_1 _5037_ (.A(_2573_),
    .Y(_2574_));
 sky130_fd_sc_hs__inv_1 _5038_ (.A(_2596_),
    .Y(_2604_));
 sky130_fd_sc_hs__inv_1 _5039_ (.A(_2601_),
    .Y(_2602_));
 sky130_fd_sc_hs__inv_1 _5040_ (.A(_2611_),
    .Y(_2613_));
 sky130_fd_sc_hs__inv_1 _5041_ (.A(_2623_),
    .Y(_2631_));
 sky130_fd_sc_hs__inv_1 _5042_ (.A(_2628_),
    .Y(_2629_));
 sky130_fd_sc_hs__inv_1 _5043_ (.A(_2654_),
    .Y(_2662_));
 sky130_fd_sc_hs__inv_1 _5044_ (.A(_2659_),
    .Y(_2660_));
 sky130_fd_sc_hs__inv_1 _5045_ (.A(_2669_),
    .Y(_2671_));
 sky130_fd_sc_hs__inv_1 _5046_ (.A(_2681_),
    .Y(_2689_));
 sky130_fd_sc_hs__inv_1 _5047_ (.A(_2686_),
    .Y(_2687_));
 sky130_fd_sc_hs__inv_1 _5048_ (.A(_2707_),
    .Y(_2715_));
 sky130_fd_sc_hs__inv_1 _5049_ (.A(_2712_),
    .Y(_2713_));
 sky130_fd_sc_hs__inv_1 _5050_ (.A(_2722_),
    .Y(_2724_));
 sky130_fd_sc_hs__inv_1 _5051_ (.A(_2734_),
    .Y(_2742_));
 sky130_fd_sc_hs__inv_1 _5052_ (.A(_2739_),
    .Y(_2740_));
 sky130_fd_sc_hs__inv_1 _5053_ (.A(_2756_),
    .Y(_2759_));
 sky130_fd_sc_hs__inv_1 _5054_ (.A(_2766_),
    .Y(_2767_));
 sky130_fd_sc_hs__inv_1 _5055_ (.A(_2777_),
    .Y(_2787_));
 sky130_fd_sc_hs__inv_1 _5056_ (.A(_2784_),
    .Y(_2785_));
 sky130_fd_sc_hs__inv_1 _5057_ (.A(_2794_),
    .Y(_2796_));
 sky130_fd_sc_hs__inv_1 _5058_ (.A(_2806_),
    .Y(_2814_));
 sky130_fd_sc_hs__inv_1 _5059_ (.A(_2811_),
    .Y(_2812_));
 sky130_fd_sc_hs__inv_1 _5060_ (.A(_2825_),
    .Y(_2827_));
 sky130_fd_sc_hs__inv_1 _5061_ (.A(_2841_),
    .Y(_2849_));
 sky130_fd_sc_hs__inv_1 _5062_ (.A(_2846_),
    .Y(_2847_));
 sky130_fd_sc_hs__inv_1 _5063_ (.A(_2856_),
    .Y(_2858_));
 sky130_fd_sc_hs__inv_1 _5064_ (.A(_2868_),
    .Y(_2876_));
 sky130_fd_sc_hs__inv_1 _5065_ (.A(_2873_),
    .Y(_2874_));
 sky130_fd_sc_hs__inv_1 _5066_ (.A(_2887_),
    .Y(_2889_));
 sky130_fd_sc_hs__inv_1 _5067_ (.A(_2897_),
    .Y(_2898_));
 sky130_fd_sc_hs__inv_1 _5068_ (.A(_2905_),
    .Y(_2912_));
 sky130_fd_sc_hs__inv_1 _5069_ (.A(_2909_),
    .Y(_2910_));
 sky130_fd_sc_hs__inv_1 _5070_ (.A(_2919_),
    .Y(_2921_));
 sky130_fd_sc_hs__inv_1 _5071_ (.A(_2931_),
    .Y(_2939_));
 sky130_fd_sc_hs__inv_1 _5072_ (.A(_2936_),
    .Y(_2937_));
 sky130_fd_sc_hs__inv_1 _5073_ (.A(_2950_),
    .Y(_2952_));
 sky130_fd_sc_hs__inv_1 _5074_ (.A(_2960_),
    .Y(_2961_));
 sky130_fd_sc_hs__inv_1 _5075_ (.A(_2969_),
    .Y(_2975_));
 sky130_fd_sc_hs__inv_1 _5076_ (.A(_2982_),
    .Y(_2984_));
 sky130_fd_sc_hs__inv_1 _5077_ (.A(_2994_),
    .Y(_3002_));
 sky130_fd_sc_hs__inv_1 _5078_ (.A(_2999_),
    .Y(_3000_));
 sky130_fd_sc_hs__inv_1 _5079_ (.A(_3013_),
    .Y(_3015_));
 sky130_fd_sc_hs__inv_2 _5080_ (.A(_3023_),
    .Y(_3024_));
 sky130_fd_sc_hs__inv_1 _5081_ (.A(_3032_),
    .Y(_3034_));
 sky130_fd_sc_hs__inv_1 _5082_ (.A(_3041_),
    .Y(_3043_));
 sky130_fd_sc_hs__inv_1 _5083_ (.A(_3053_),
    .Y(_3061_));
 sky130_fd_sc_hs__inv_1 _5084_ (.A(_3058_),
    .Y(_3059_));
 sky130_fd_sc_hs__inv_1 _5085_ (.A(_3072_),
    .Y(_3074_));
 sky130_fd_sc_hs__clkinv_2 _5086_ (.A(_3082_),
    .Y(_3083_));
 sky130_fd_sc_hs__inv_1 _5087_ (.A(_3094_),
    .Y(_3103_));
 sky130_fd_sc_hs__inv_1 _5088_ (.A(_3098_),
    .Y(_3100_));
 sky130_fd_sc_hs__inv_1 _5089_ (.A(_3110_),
    .Y(_3118_));
 sky130_fd_sc_hs__inv_1 _5090_ (.A(_3115_),
    .Y(_3116_));
 sky130_fd_sc_hs__inv_1 _5091_ (.A(_3129_),
    .Y(_3131_));
 sky130_fd_sc_hs__clkinv_2 _5092_ (.A(_3139_),
    .Y(_3140_));
 sky130_fd_sc_hs__inv_1 _5093_ (.A(_3152_),
    .Y(_3161_));
 sky130_fd_sc_hs__inv_2 _5094_ (.A(_3155_),
    .Y(_3157_));
 sky130_fd_sc_hs__inv_1 _5095_ (.A(_3168_),
    .Y(_3176_));
 sky130_fd_sc_hs__inv_1 _5096_ (.A(_3173_),
    .Y(_3174_));
 sky130_fd_sc_hs__inv_1 _5097_ (.A(_3187_),
    .Y(_3189_));
 sky130_fd_sc_hs__inv_1 _5098_ (.A(_3197_),
    .Y(_3198_));
 sky130_fd_sc_hs__inv_1 _5099_ (.A(_3210_),
    .Y(_3215_));
 sky130_fd_sc_hs__inv_1 _5100_ (.A(_3222_),
    .Y(_3230_));
 sky130_fd_sc_hs__inv_1 _5101_ (.A(_3227_),
    .Y(_3228_));
 sky130_fd_sc_hs__inv_1 _5102_ (.A(_3241_),
    .Y(_3243_));
 sky130_fd_sc_hs__inv_1 _5103_ (.A(_3251_),
    .Y(_3252_));
 sky130_fd_sc_hs__inv_1 _5104_ (.A(_3267_),
    .Y(_3284_));
 sky130_fd_sc_hs__inv_1 _5105_ (.A(_3271_),
    .Y(_3279_));
 sky130_fd_sc_hs__inv_1 _5106_ (.A(_3276_),
    .Y(_3277_));
 sky130_fd_sc_hs__inv_1 _5107_ (.A(_3291_),
    .Y(_3293_));
 sky130_fd_sc_hs__inv_1 _5108_ (.A(_3301_),
    .Y(_3302_));
 sky130_fd_sc_hs__inv_1 _5109_ (.A(_3316_),
    .Y(_3333_));
 sky130_fd_sc_hs__inv_2 _5110_ (.A(_3319_),
    .Y(_3327_));
 sky130_fd_sc_hs__inv_1 _5111_ (.A(_3324_),
    .Y(_3325_));
 sky130_fd_sc_hs__inv_1 _5112_ (.A(_3340_),
    .Y(_3342_));
 sky130_fd_sc_hs__inv_1 _5113_ (.A(_3350_),
    .Y(_3351_));
 sky130_fd_sc_hs__inv_1 _5114_ (.A(_3369_),
    .Y(_3370_));
 sky130_fd_sc_hs__inv_1 _5115_ (.A(_3383_),
    .Y(_3385_));
 sky130_fd_sc_hs__inv_1 _5116_ (.A(_3393_),
    .Y(_3394_));
 sky130_fd_sc_hs__inv_1 _5117_ (.A(_3410_),
    .Y(_3411_));
 sky130_fd_sc_hs__inv_1 _5118_ (.A(_3422_),
    .Y(_3424_));
 sky130_fd_sc_hs__inv_1 _5119_ (.A(_3432_),
    .Y(_3433_));
 sky130_fd_sc_hs__inv_1 _5120_ (.A(_3448_),
    .Y(_3449_));
 sky130_fd_sc_hs__inv_1 _5121_ (.A(_3460_),
    .Y(_3462_));
 sky130_fd_sc_hs__inv_1 _5122_ (.A(_3470_),
    .Y(_3471_));
 sky130_fd_sc_hs__inv_1 _5123_ (.A(_3490_),
    .Y(_3507_));
 sky130_fd_sc_hs__inv_1 _5124_ (.A(_3495_),
    .Y(_3497_));
 sky130_fd_sc_hs__inv_1 _5125_ (.A(_3505_),
    .Y(_3506_));
 sky130_fd_sc_hs__inv_1 _5126_ (.A(_3525_),
    .Y(_3527_));
 sky130_fd_sc_hs__inv_1 _5127_ (.A(_3534_),
    .Y(_3535_));
 sky130_fd_sc_hs__inv_1 _5128_ (.A(_3559_),
    .Y(_3560_));
 sky130_fd_sc_hs__inv_1 _5129_ (.A(_2248_),
    .Y(_2265_));
 sky130_fd_sc_hs__inv_1 _5130_ (.A(_2257_),
    .Y(_2284_));
 sky130_fd_sc_hs__inv_1 _5131_ (.A(_2277_),
    .Y(_2302_));
 sky130_fd_sc_hs__inv_1 _5132_ (.A(_2282_),
    .Y(_3743_));
 sky130_fd_sc_hs__inv_1 _5133_ (.A(_2294_),
    .Y(_2324_));
 sky130_fd_sc_hs__inv_1 _5134_ (.A(_2316_),
    .Y(_2359_));
 sky130_fd_sc_hs__inv_1 _5135_ (.A(_2351_),
    .Y(_2387_));
 sky130_fd_sc_hs__inv_1 _5136_ (.A(_2379_),
    .Y(_2419_));
 sky130_fd_sc_hs__inv_1 _5137_ (.A(_2384_),
    .Y(_2430_));
 sky130_fd_sc_hs__inv_1 _5138_ (.A(_2394_),
    .Y(_2428_));
 sky130_fd_sc_hs__inv_1 _5139_ (.A(_2411_),
    .Y(_2457_));
 sky130_fd_sc_hs__inv_1 _5140_ (.A(_2416_),
    .Y(_2468_));
 sky130_fd_sc_hs__inv_1 _5141_ (.A(_2426_),
    .Y(_2466_));
 sky130_fd_sc_hs__inv_1 _5142_ (.A(_2449_),
    .Y(_2502_));
 sky130_fd_sc_hs__inv_1 _5143_ (.A(_2454_),
    .Y(_2513_));
 sky130_fd_sc_hs__inv_1 _5144_ (.A(_2464_),
    .Y(_2511_));
 sky130_fd_sc_hs__inv_1 _5145_ (.A(_2476_),
    .Y(_2524_));
 sky130_fd_sc_hs__inv_1 _5146_ (.A(_2479_),
    .Y(_2528_));
 sky130_fd_sc_hs__inv_1 _5147_ (.A(_2494_),
    .Y(_2548_));
 sky130_fd_sc_hs__inv_1 _5148_ (.A(_2499_),
    .Y(_2559_));
 sky130_fd_sc_hs__inv_1 _5149_ (.A(_2509_),
    .Y(_2557_));
 sky130_fd_sc_hs__inv_1 _5150_ (.A(_2521_),
    .Y(_2575_));
 sky130_fd_sc_hs__inv_1 _5151_ (.A(_2540_),
    .Y(_2603_));
 sky130_fd_sc_hs__inv_1 _5152_ (.A(_2545_),
    .Y(_2614_));
 sky130_fd_sc_hs__inv_1 _5153_ (.A(_2555_),
    .Y(_2612_));
 sky130_fd_sc_hs__inv_1 _5154_ (.A(_2567_),
    .Y(_2630_));
 sky130_fd_sc_hs__inv_1 _5155_ (.A(_2590_),
    .Y(_2646_));
 sky130_fd_sc_hs__inv_1 _5156_ (.A(_2595_),
    .Y(_2661_));
 sky130_fd_sc_hs__inv_1 _5157_ (.A(_2600_),
    .Y(_2672_));
 sky130_fd_sc_hs__inv_1 _5158_ (.A(_2610_),
    .Y(_2670_));
 sky130_fd_sc_hs__inv_1 _5159_ (.A(_2622_),
    .Y(_2688_));
 sky130_fd_sc_hs__inv_1 _5160_ (.A(_2653_),
    .Y(_2714_));
 sky130_fd_sc_hs__inv_1 _5161_ (.A(_2658_),
    .Y(_2725_));
 sky130_fd_sc_hs__inv_1 _5162_ (.A(_2668_),
    .Y(_2723_));
 sky130_fd_sc_hs__inv_1 _5163_ (.A(_2680_),
    .Y(_2741_));
 sky130_fd_sc_hs__inv_1 _5164_ (.A(_2706_),
    .Y(_2786_));
 sky130_fd_sc_hs__inv_1 _5165_ (.A(_2711_),
    .Y(_2797_));
 sky130_fd_sc_hs__inv_1 _5166_ (.A(_2721_),
    .Y(_2795_));
 sky130_fd_sc_hs__inv_1 _5167_ (.A(_2733_),
    .Y(_2813_));
 sky130_fd_sc_hs__inv_1 _5168_ (.A(_2738_),
    .Y(_2828_));
 sky130_fd_sc_hs__inv_1 _5169_ (.A(_2752_),
    .Y(_2826_));
 sky130_fd_sc_hs__inv_1 _5170_ (.A(_2765_),
    .Y(_2836_));
 sky130_fd_sc_hs__inv_1 _5171_ (.A(_2776_),
    .Y(_2848_));
 sky130_fd_sc_hs__inv_1 _5172_ (.A(_2783_),
    .Y(_2859_));
 sky130_fd_sc_hs__inv_1 _5173_ (.A(_2793_),
    .Y(_2857_));
 sky130_fd_sc_hs__inv_1 _5174_ (.A(_2805_),
    .Y(_2875_));
 sky130_fd_sc_hs__inv_1 _5175_ (.A(_2810_),
    .Y(_2890_));
 sky130_fd_sc_hs__inv_1 _5176_ (.A(_2824_),
    .Y(_2888_));
 sky130_fd_sc_hs__inv_1 _5177_ (.A(_2840_),
    .Y(_2911_));
 sky130_fd_sc_hs__inv_1 _5178_ (.A(_2845_),
    .Y(_2922_));
 sky130_fd_sc_hs__inv_1 _5179_ (.A(_2855_),
    .Y(_2920_));
 sky130_fd_sc_hs__inv_1 _5180_ (.A(_2867_),
    .Y(_2938_));
 sky130_fd_sc_hs__inv_1 _5181_ (.A(_2872_),
    .Y(_2953_));
 sky130_fd_sc_hs__inv_1 _5182_ (.A(_2886_),
    .Y(_2951_));
 sky130_fd_sc_hs__inv_1 _5183_ (.A(_2896_),
    .Y(_2964_));
 sky130_fd_sc_hs__inv_1 _5184_ (.A(_2904_),
    .Y(_2974_));
 sky130_fd_sc_hs__inv_1 _5185_ (.A(_2908_),
    .Y(_2985_));
 sky130_fd_sc_hs__inv_1 _5186_ (.A(_2918_),
    .Y(_2983_));
 sky130_fd_sc_hs__inv_1 _5187_ (.A(_2930_),
    .Y(_3001_));
 sky130_fd_sc_hs__inv_1 _5188_ (.A(_2935_),
    .Y(_3016_));
 sky130_fd_sc_hs__inv_1 _5189_ (.A(_2949_),
    .Y(_3014_));
 sky130_fd_sc_hs__clkinv_2 _5190_ (.A(_2959_),
    .Y(_3027_));
 sky130_fd_sc_hs__inv_1 _5191_ (.A(_2968_),
    .Y(_3033_));
 sky130_fd_sc_hs__inv_2 _5192_ (.A(_2971_),
    .Y(_3044_));
 sky130_fd_sc_hs__inv_1 _5193_ (.A(_2981_),
    .Y(_3042_));
 sky130_fd_sc_hs__inv_1 _5194_ (.A(_2993_),
    .Y(_3060_));
 sky130_fd_sc_hs__inv_1 _5195_ (.A(_2998_),
    .Y(_3075_));
 sky130_fd_sc_hs__inv_1 _5196_ (.A(_3012_),
    .Y(_3073_));
 sky130_fd_sc_hs__clkinv_2 _5197_ (.A(_3022_),
    .Y(_3086_));
 sky130_fd_sc_hs__inv_1 _5198_ (.A(_3040_),
    .Y(_3099_));
 sky130_fd_sc_hs__inv_1 _5199_ (.A(_3052_),
    .Y(_3117_));
 sky130_fd_sc_hs__inv_1 _5200_ (.A(_3057_),
    .Y(_3132_));
 sky130_fd_sc_hs__inv_1 _5201_ (.A(_3071_),
    .Y(_3130_));
 sky130_fd_sc_hs__inv_2 _5202_ (.A(_3081_),
    .Y(_3143_));
 sky130_fd_sc_hs__inv_1 _5203_ (.A(_3093_),
    .Y(_3160_));
 sky130_fd_sc_hs__inv_1 _5204_ (.A(_3097_),
    .Y(_3156_));
 sky130_fd_sc_hs__inv_1 _5205_ (.A(_3109_),
    .Y(_3175_));
 sky130_fd_sc_hs__inv_1 _5206_ (.A(_3114_),
    .Y(_3190_));
 sky130_fd_sc_hs__inv_1 _5207_ (.A(_3128_),
    .Y(_3188_));
 sky130_fd_sc_hs__inv_1 _5208_ (.A(_3138_),
    .Y(_3201_));
 sky130_fd_sc_hs__inv_1 _5209_ (.A(_3151_),
    .Y(_3214_));
 sky130_fd_sc_hs__inv_1 _5210_ (.A(_3154_),
    .Y(_3211_));
 sky130_fd_sc_hs__inv_1 _5211_ (.A(_3167_),
    .Y(_3229_));
 sky130_fd_sc_hs__inv_1 _5212_ (.A(_3172_),
    .Y(_3244_));
 sky130_fd_sc_hs__inv_1 _5213_ (.A(_3186_),
    .Y(_3242_));
 sky130_fd_sc_hs__clkinv_2 _5214_ (.A(_3196_),
    .Y(_3255_));
 sky130_fd_sc_hs__inv_1 _5215_ (.A(_3221_),
    .Y(_3278_));
 sky130_fd_sc_hs__inv_1 _5216_ (.A(_3226_),
    .Y(_3294_));
 sky130_fd_sc_hs__inv_1 _5217_ (.A(_3240_),
    .Y(_3292_));
 sky130_fd_sc_hs__inv_1 _5218_ (.A(_3250_),
    .Y(_3305_));
 sky130_fd_sc_hs__inv_1 _5219_ (.A(_3266_),
    .Y(_3332_));
 sky130_fd_sc_hs__inv_1 _5220_ (.A(_3270_),
    .Y(_3326_));
 sky130_fd_sc_hs__inv_1 _5221_ (.A(_3275_),
    .Y(_3343_));
 sky130_fd_sc_hs__inv_1 _5222_ (.A(_3290_),
    .Y(_3341_));
 sky130_fd_sc_hs__inv_1 _5223_ (.A(_3300_),
    .Y(_3354_));
 sky130_fd_sc_hs__inv_1 _5224_ (.A(_3312_),
    .Y(_3362_));
 sky130_fd_sc_hs__inv_1 _5225_ (.A(_3315_),
    .Y(_3376_));
 sky130_fd_sc_hs__inv_2 _5226_ (.A(_3318_),
    .Y(_3371_));
 sky130_fd_sc_hs__inv_1 _5227_ (.A(_3323_),
    .Y(_3386_));
 sky130_fd_sc_hs__inv_1 _5228_ (.A(_3339_),
    .Y(_3384_));
 sky130_fd_sc_hs__inv_1 _5229_ (.A(_3349_),
    .Y(_3397_));
 sky130_fd_sc_hs__inv_1 _5230_ (.A(_3368_),
    .Y(_3425_));
 sky130_fd_sc_hs__inv_1 _5231_ (.A(_3382_),
    .Y(_3423_));
 sky130_fd_sc_hs__inv_1 _5232_ (.A(_3392_),
    .Y(_3436_));
 sky130_fd_sc_hs__inv_1 _5233_ (.A(_3409_),
    .Y(_3463_));
 sky130_fd_sc_hs__inv_1 _5234_ (.A(_3421_),
    .Y(_3461_));
 sky130_fd_sc_hs__inv_1 _5235_ (.A(_3431_),
    .Y(_3474_));
 sky130_fd_sc_hs__inv_1 _5236_ (.A(_3447_),
    .Y(_3498_));
 sky130_fd_sc_hs__inv_1 _5237_ (.A(_3459_),
    .Y(_3496_));
 sky130_fd_sc_hs__inv_1 _5238_ (.A(_3469_),
    .Y(_3510_));
 sky130_fd_sc_hs__inv_1 _5239_ (.A(_3489_),
    .Y(_3536_));
 sky130_fd_sc_hs__inv_1 _5240_ (.A(_3494_),
    .Y(_3526_));
 sky130_fd_sc_hs__inv_1 _5241_ (.A(_3504_),
    .Y(_3539_));
 sky130_fd_sc_hs__inv_1 _5242_ (.A(_3533_),
    .Y(_3563_));
 sky130_fd_sc_hs__inv_1 _5243_ (.A(net74),
    .Y(_3566_));
 sky130_fd_sc_hs__clkbuf_4 _5244_ (.A(_0107_),
    .X(_0568_));
 sky130_fd_sc_hs__nor2_4 _5245_ (.A(_0106_),
    .B(_0387_),
    .Y(_0569_));
 sky130_fd_sc_hs__clkbuf_4 _5246_ (.A(_0569_),
    .X(_0570_));
 sky130_fd_sc_hs__a22o_2 _5247_ (.A1(net2),
    .A2(_0568_),
    .B1(_0570_),
    .B2(_0435_),
    .X(_2227_));
 sky130_fd_sc_hs__a22o_1 _5248_ (.A1(net21),
    .A2(_0568_),
    .B1(_0570_),
    .B2(_0447_),
    .X(_3578_));
 sky130_fd_sc_hs__a22o_1 _5249_ (.A1(net32),
    .A2(_0568_),
    .B1(_0570_),
    .B2(_0450_),
    .X(_3582_));
 sky130_fd_sc_hs__clkbuf_4 _5250_ (.A(_0107_),
    .X(_0571_));
 sky130_fd_sc_hs__buf_8 _5251_ (.A(imd_val_q_i[37]),
    .X(_0572_));
 sky130_fd_sc_hs__a22o_1 _5252_ (.A1(net35),
    .A2(_0571_),
    .B1(_0570_),
    .B2(_0572_),
    .X(_3586_));
 sky130_fd_sc_hs__buf_8 _5253_ (.A(imd_val_q_i[38]),
    .X(_0573_));
 sky130_fd_sc_hs__a22o_1 _5254_ (.A1(net36),
    .A2(_0571_),
    .B1(_0570_),
    .B2(_0573_),
    .X(_3590_));
 sky130_fd_sc_hs__clkbuf_16 _5255_ (.A(imd_val_q_i[39]),
    .X(_0574_));
 sky130_fd_sc_hs__a22o_1 _5256_ (.A1(net37),
    .A2(_0571_),
    .B1(_0570_),
    .B2(_0574_),
    .X(_3594_));
 sky130_fd_sc_hs__clkbuf_16 _5257_ (.A(imd_val_q_i[40]),
    .X(_0575_));
 sky130_fd_sc_hs__a22o_2 _5258_ (.A1(net38),
    .A2(_0571_),
    .B1(_0570_),
    .B2(_0575_),
    .X(_3598_));
 sky130_fd_sc_hs__clkbuf_16 _5259_ (.A(imd_val_q_i[41]),
    .X(_0576_));
 sky130_fd_sc_hs__a22o_4 _5260_ (.A1(net39),
    .A2(_0571_),
    .B1(_0570_),
    .B2(_0576_),
    .X(_3602_));
 sky130_fd_sc_hs__clkbuf_16 _5261_ (.A(imd_val_q_i[42]),
    .X(_0577_));
 sky130_fd_sc_hs__a22o_2 _5262_ (.A1(net40),
    .A2(_0571_),
    .B1(_0570_),
    .B2(_0577_),
    .X(_3606_));
 sky130_fd_sc_hs__buf_8 _5263_ (.A(imd_val_q_i[43]),
    .X(_0578_));
 sky130_fd_sc_hs__a22o_1 _5264_ (.A1(net41),
    .A2(_0571_),
    .B1(_0570_),
    .B2(_0578_),
    .X(_3610_));
 sky130_fd_sc_hs__clkbuf_4 _5265_ (.A(_0569_),
    .X(_0579_));
 sky130_fd_sc_hs__clkbuf_16 _5266_ (.A(imd_val_q_i[44]),
    .X(_0580_));
 sky130_fd_sc_hs__a22o_1 _5267_ (.A1(net3),
    .A2(_0571_),
    .B1(_0579_),
    .B2(_0580_),
    .X(_3614_));
 sky130_fd_sc_hs__buf_16 _5268_ (.A(imd_val_q_i[45]),
    .X(_0581_));
 sky130_fd_sc_hs__a22o_2 _5269_ (.A1(net4),
    .A2(_0571_),
    .B1(_0579_),
    .B2(_0581_),
    .X(_3618_));
 sky130_fd_sc_hs__buf_16 _5270_ (.A(imd_val_q_i[46]),
    .X(_0582_));
 sky130_fd_sc_hs__a22o_2 _5271_ (.A1(net5),
    .A2(_0571_),
    .B1(_0579_),
    .B2(_0582_),
    .X(_3622_));
 sky130_fd_sc_hs__clkbuf_4 _5272_ (.A(_0106_),
    .X(_0583_));
 sky130_fd_sc_hs__clkbuf_16 _5273_ (.A(imd_val_q_i[47]),
    .X(_0584_));
 sky130_fd_sc_hs__a22o_2 _5274_ (.A1(net6),
    .A2(_0583_),
    .B1(_0579_),
    .B2(_0584_),
    .X(_3626_));
 sky130_fd_sc_hs__buf_8 _5275_ (.A(imd_val_q_i[48]),
    .X(_0585_));
 sky130_fd_sc_hs__a22o_2 _5276_ (.A1(net7),
    .A2(_0583_),
    .B1(_0579_),
    .B2(_0585_),
    .X(_3630_));
 sky130_fd_sc_hs__a22o_2 _5277_ (.A1(net8),
    .A2(_0583_),
    .B1(_0579_),
    .B2(net107),
    .X(_3634_));
 sky130_fd_sc_hs__a22o_2 _5278_ (.A1(net17),
    .A2(_0583_),
    .B1(_0579_),
    .B2(_0436_),
    .X(_3638_));
 sky130_fd_sc_hs__a22o_2 _5279_ (.A1(net18),
    .A2(_0583_),
    .B1(_0579_),
    .B2(_0446_),
    .X(_3642_));
 sky130_fd_sc_hs__a22o_1 _5280_ (.A1(net19),
    .A2(_0583_),
    .B1(_0579_),
    .B2(_0449_),
    .X(_3646_));
 sky130_fd_sc_hs__clkbuf_16 _5281_ (.A(imd_val_q_i[53]),
    .X(_0586_));
 sky130_fd_sc_hs__a22o_1 _5282_ (.A1(net20),
    .A2(_0583_),
    .B1(_0579_),
    .B2(_0586_),
    .X(_3650_));
 sky130_fd_sc_hs__clkbuf_4 _5283_ (.A(_0569_),
    .X(_0587_));
 sky130_fd_sc_hs__clkbuf_16 _5284_ (.A(imd_val_q_i[54]),
    .X(_0588_));
 sky130_fd_sc_hs__a22o_2 _5285_ (.A1(net22),
    .A2(_0583_),
    .B1(_0587_),
    .B2(_0588_),
    .X(_3654_));
 sky130_fd_sc_hs__a22o_2 _5286_ (.A1(net23),
    .A2(_0583_),
    .B1(_0587_),
    .B2(net109),
    .X(_3658_));
 sky130_fd_sc_hs__a22o_1 _5287_ (.A1(net24),
    .A2(_0583_),
    .B1(_0587_),
    .B2(_0520_),
    .X(_3662_));
 sky130_fd_sc_hs__a22o_1 _5288_ (.A1(net25),
    .A2(_0108_),
    .B1(_0587_),
    .B2(_0526_),
    .X(_3666_));
 sky130_fd_sc_hs__a22o_1 _5289_ (.A1(net26),
    .A2(_0108_),
    .B1(_0587_),
    .B2(_0527_),
    .X(_3670_));
 sky130_fd_sc_hs__a22o_1 _5290_ (.A1(net27),
    .A2(_0108_),
    .B1(_0587_),
    .B2(_0529_),
    .X(_3674_));
 sky130_fd_sc_hs__a22o_1 _5291_ (.A1(net28),
    .A2(_0108_),
    .B1(_0587_),
    .B2(_0565_),
    .X(_3678_));
 sky130_fd_sc_hs__a22o_1 _5292_ (.A1(net29),
    .A2(_0108_),
    .B1(_0587_),
    .B2(_0566_),
    .X(_3682_));
 sky130_fd_sc_hs__a22o_1 _5293_ (.A1(net30),
    .A2(_0108_),
    .B1(_0587_),
    .B2(net111),
    .X(_3686_));
 sky130_fd_sc_hs__a22o_1 _5294_ (.A1(net31),
    .A2(_0108_),
    .B1(_0587_),
    .B2(net112),
    .X(_3690_));
 sky130_fd_sc_hs__a22o_1 _5295_ (.A1(net33),
    .A2(_0108_),
    .B1(_0569_),
    .B2(_0567_),
    .X(_3694_));
 sky130_fd_sc_hs__clkbuf_4 _5296_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .X(_0589_));
 sky130_fd_sc_hs__buf_8 _5297_ (.A(_0589_),
    .X(_0590_));
 sky130_fd_sc_hs__inv_2 _5298_ (.A(_0590_),
    .Y(_3702_));
 sky130_fd_sc_hs__inv_1 _5299_ (.A(_2233_),
    .Y(_2241_));
 sky130_fd_sc_hs__inv_1 _5300_ (.A(_2252_),
    .Y(_2270_));
 sky130_fd_sc_hs__inv_1 _5301_ (.A(_2310_),
    .Y(_3750_));
 sky130_fd_sc_hs__inv_1 _5302_ (.A(_2340_),
    .Y(_3759_));
 sky130_fd_sc_hs__nor2_1 _5303_ (.A(_0460_),
    .B(_0482_),
    .Y(_2376_));
 sky130_fd_sc_hs__nor2_1 _5304_ (.A(_0460_),
    .B(_0486_),
    .Y(_2408_));
 sky130_fd_sc_hs__inv_1 _5305_ (.A(_2405_),
    .Y(_3781_));
 sky130_fd_sc_hs__nor2_1 _5306_ (.A(_0460_),
    .B(_0490_),
    .Y(_2446_));
 sky130_fd_sc_hs__inv_1 _5307_ (.A(_2444_),
    .Y(_3787_));
 sky130_fd_sc_hs__nor2_2 _5308_ (.A(_0459_),
    .B(_0493_),
    .Y(_2491_));
 sky130_fd_sc_hs__inv_1 _5309_ (.A(_2486_),
    .Y(_2533_));
 sky130_fd_sc_hs__inv_1 _5310_ (.A(_2489_),
    .Y(_3797_));
 sky130_fd_sc_hs__nor2_2 _5311_ (.A(_0459_),
    .B(_0497_),
    .Y(_2537_));
 sky130_fd_sc_hs__inv_1 _5312_ (.A(_2578_),
    .Y(_2580_));
 sky130_fd_sc_hs__inv_1 _5313_ (.A(_2526_),
    .Y(_2579_));
 sky130_fd_sc_hs__inv_1 _5314_ (.A(_2531_),
    .Y(_2588_));
 sky130_fd_sc_hs__nor2_2 _5315_ (.A(_0459_),
    .B(_0501_),
    .Y(_2592_));
 sky130_fd_sc_hs__inv_1 _5316_ (.A(_2633_),
    .Y(_2635_));
 sky130_fd_sc_hs__inv_1 _5317_ (.A(_2577_),
    .Y(_2634_));
 sky130_fd_sc_hs__nor2_2 _5318_ (.A(_0459_),
    .B(_0505_),
    .Y(_2650_));
 sky130_fd_sc_hs__inv_1 _5319_ (.A(_2647_),
    .Y(_3821_));
 sky130_fd_sc_hs__inv_1 _5320_ (.A(_2761_),
    .Y(_2763_));
 sky130_fd_sc_hs__inv_1 _5321_ (.A(_2700_),
    .Y(_3825_));
 sky130_fd_sc_hs__inv_1 _5322_ (.A(_2771_),
    .Y(_3831_));
 sky130_fd_sc_hs__nand2_1 _5323_ (.A(_0449_),
    .B(_0086_),
    .Y(_0591_));
 sky130_fd_sc_hs__nand2_4 _5324_ (.A(_0528_),
    .B(_0591_),
    .Y(_2839_));
 sky130_fd_sc_hs__inv_1 _5325_ (.A(_2829_),
    .Y(_3835_));
 sky130_fd_sc_hs__inv_1 _5326_ (.A(_2837_),
    .Y(_3837_));
 sky130_fd_sc_hs__nand2_1 _5327_ (.A(_0586_),
    .B(_0086_),
    .Y(_0592_));
 sky130_fd_sc_hs__nand2_2 _5328_ (.A(_0528_),
    .B(_0592_),
    .Y(_2903_));
 sky130_fd_sc_hs__inv_1 _5329_ (.A(_2891_),
    .Y(_3841_));
 sky130_fd_sc_hs__inv_1 _5330_ (.A(_2901_),
    .Y(_3843_));
 sky130_fd_sc_hs__nand2_1 _5331_ (.A(_0588_),
    .B(_0086_),
    .Y(_0593_));
 sky130_fd_sc_hs__nand2_2 _5332_ (.A(_0528_),
    .B(_0593_),
    .Y(_2967_));
 sky130_fd_sc_hs__inv_1 _5333_ (.A(_2954_),
    .Y(_3847_));
 sky130_fd_sc_hs__inv_1 _5334_ (.A(_2965_),
    .Y(_3849_));
 sky130_fd_sc_hs__nand2_1 _5335_ (.A(net109),
    .B(_0086_),
    .Y(_0594_));
 sky130_fd_sc_hs__nand2_2 _5336_ (.A(_0528_),
    .B(_0594_),
    .Y(_3030_));
 sky130_fd_sc_hs__inv_1 _5337_ (.A(_3017_),
    .Y(_3853_));
 sky130_fd_sc_hs__inv_1 _5338_ (.A(_3028_),
    .Y(_3855_));
 sky130_fd_sc_hs__inv_1 _5339_ (.A(_3076_),
    .Y(_3859_));
 sky130_fd_sc_hs__inv_1 _5340_ (.A(_3087_),
    .Y(_3861_));
 sky130_fd_sc_hs__inv_1 _5341_ (.A(_3090_),
    .Y(_3149_));
 sky130_fd_sc_hs__inv_1 _5342_ (.A(_3133_),
    .Y(_3865_));
 sky130_fd_sc_hs__inv_1 _5343_ (.A(_3144_),
    .Y(_3867_));
 sky130_fd_sc_hs__inv_1 _5344_ (.A(_3147_),
    .Y(_3207_));
 sky130_fd_sc_hs__inv_1 _5345_ (.A(_3191_),
    .Y(_3871_));
 sky130_fd_sc_hs__inv_1 _5346_ (.A(_3202_),
    .Y(_3873_));
 sky130_fd_sc_hs__inv_1 _5347_ (.A(_3245_),
    .Y(_3877_));
 sky130_fd_sc_hs__inv_1 _5348_ (.A(_3256_),
    .Y(_3879_));
 sky130_fd_sc_hs__inv_1 _5349_ (.A(_3262_),
    .Y(_3314_));
 sky130_fd_sc_hs__inv_1 _5350_ (.A(_3295_),
    .Y(_3883_));
 sky130_fd_sc_hs__inv_1 _5351_ (.A(_3306_),
    .Y(_3885_));
 sky130_fd_sc_hs__inv_1 _5352_ (.A(_3344_),
    .Y(_3889_));
 sky130_fd_sc_hs__inv_1 _5353_ (.A(_3355_),
    .Y(_3891_));
 sky130_fd_sc_hs__inv_1 _5354_ (.A(_3387_),
    .Y(_3895_));
 sky130_fd_sc_hs__inv_1 _5355_ (.A(_3398_),
    .Y(_3897_));
 sky130_fd_sc_hs__inv_1 _5356_ (.A(_3426_),
    .Y(_3901_));
 sky130_fd_sc_hs__inv_1 _5357_ (.A(_3437_),
    .Y(_3903_));
 sky130_fd_sc_hs__inv_1 _5358_ (.A(_3444_),
    .Y(_3487_));
 sky130_fd_sc_hs__inv_1 _5359_ (.A(_3464_),
    .Y(_3907_));
 sky130_fd_sc_hs__inv_1 _5360_ (.A(_3475_),
    .Y(_3909_));
 sky130_fd_sc_hs__inv_1 _5361_ (.A(_3499_),
    .Y(_3913_));
 sky130_fd_sc_hs__inv_1 _5362_ (.A(_3511_),
    .Y(_3915_));
 sky130_fd_sc_hs__inv_1 _5363_ (.A(_3528_),
    .Y(_3921_));
 sky130_fd_sc_hs__inv_1 _5364_ (.A(_3540_),
    .Y(_3923_));
 sky130_fd_sc_hs__inv_1 _5365_ (.A(net75),
    .Y(_3567_));
 sky130_fd_sc_hs__clkbuf_16 _5366_ (.A(_0107_),
    .X(_0595_));
 sky130_fd_sc_hs__buf_8 _5367_ (.A(_0561_),
    .X(_0596_));
 sky130_fd_sc_hs__nand2_8 _5368_ (.A(_0116_),
    .B(_0121_),
    .Y(_0597_));
 sky130_fd_sc_hs__buf_16 _5369_ (.A(_0597_),
    .X(_0598_));
 sky130_fd_sc_hs__xnor2_2 _5370_ (.A(_0596_),
    .B(_0598_),
    .Y(_0599_));
 sky130_fd_sc_hs__clkbuf_16 _5371_ (.A(_0107_),
    .X(_0600_));
 sky130_fd_sc_hs__buf_8 _5372_ (.A(net366),
    .X(_0601_));
 sky130_fd_sc_hs__clkbuf_8 _5373_ (.A(net366),
    .X(_0602_));
 sky130_fd_sc_hs__buf_4 _5374_ (.A(_0387_),
    .X(_0603_));
 sky130_fd_sc_hs__nor2_1 _5375_ (.A(net81),
    .B(_0603_),
    .Y(_0604_));
 sky130_fd_sc_hs__clkbuf_16 _5376_ (.A(_0381_),
    .X(_0605_));
 sky130_fd_sc_hs__o22ai_4 _5377_ (.A1(_0605_),
    .A2(_0435_),
    .B1(net121),
    .B2(_0427_),
    .Y(_0606_));
 sky130_fd_sc_hs__nor3_2 _5378_ (.A(_0602_),
    .B(_0604_),
    .C(_0606_),
    .Y(_0607_));
 sky130_fd_sc_hs__a21oi_4 _5379_ (.A1(net153),
    .A2(_0601_),
    .B1(_0607_),
    .Y(_0608_));
 sky130_fd_sc_hs__nor2_8 _5380_ (.A(_0600_),
    .B(_0608_),
    .Y(_0609_));
 sky130_fd_sc_hs__a21oi_4 _5381_ (.A1(_0595_),
    .A2(_0599_),
    .B1(_0609_),
    .Y(_2228_));
 sky130_fd_sc_hs__xnor2_1 _5382_ (.A(net53),
    .B(_0598_),
    .Y(_0610_));
 sky130_fd_sc_hs__nor2_1 _5383_ (.A(net92),
    .B(_0603_),
    .Y(_0611_));
 sky130_fd_sc_hs__o22ai_4 _5384_ (.A1(_0605_),
    .A2(_0447_),
    .B1(net132),
    .B2(_0427_),
    .Y(_0612_));
 sky130_fd_sc_hs__nor3_1 _5385_ (.A(_0602_),
    .B(_0611_),
    .C(_0612_),
    .Y(_0613_));
 sky130_fd_sc_hs__a21oi_2 _5386_ (.A1(net164),
    .A2(_0601_),
    .B1(_0613_),
    .Y(_0614_));
 sky130_fd_sc_hs__nor2_4 _5387_ (.A(_0600_),
    .B(_0614_),
    .Y(_0615_));
 sky130_fd_sc_hs__a21oi_1 _5388_ (.A1(_0595_),
    .A2(_0610_),
    .B1(_0615_),
    .Y(_3579_));
 sky130_fd_sc_hs__xnor2_1 _5389_ (.A(net64),
    .B(_0598_),
    .Y(_0616_));
 sky130_fd_sc_hs__nor2_1 _5390_ (.A(net103),
    .B(_0603_),
    .Y(_0617_));
 sky130_fd_sc_hs__o22ai_2 _5391_ (.A1(_0605_),
    .A2(_0450_),
    .B1(net143),
    .B2(_0427_),
    .Y(_0618_));
 sky130_fd_sc_hs__nor3_2 _5392_ (.A(_0602_),
    .B(_0617_),
    .C(_0618_),
    .Y(_0619_));
 sky130_fd_sc_hs__a21oi_4 _5393_ (.A1(net175),
    .A2(_0601_),
    .B1(_0619_),
    .Y(_0620_));
 sky130_fd_sc_hs__nor2_4 _5394_ (.A(_0600_),
    .B(_0620_),
    .Y(_0621_));
 sky130_fd_sc_hs__a21oi_1 _5395_ (.A1(_0595_),
    .A2(_0616_),
    .B1(_0621_),
    .Y(_3583_));
 sky130_fd_sc_hs__xnor2_2 _5396_ (.A(net67),
    .B(_0598_),
    .Y(_0622_));
 sky130_fd_sc_hs__nor2_1 _5397_ (.A(net106),
    .B(_0603_),
    .Y(_0623_));
 sky130_fd_sc_hs__o22ai_4 _5398_ (.A1(_0605_),
    .A2(_0572_),
    .B1(net146),
    .B2(_0427_),
    .Y(_0624_));
 sky130_fd_sc_hs__nor3_1 _5399_ (.A(_0602_),
    .B(_0623_),
    .C(_0624_),
    .Y(_0625_));
 sky130_fd_sc_hs__a21oi_2 _5400_ (.A1(net178),
    .A2(_0601_),
    .B1(_0625_),
    .Y(_0626_));
 sky130_fd_sc_hs__nor2_4 _5401_ (.A(_0600_),
    .B(_0626_),
    .Y(_0627_));
 sky130_fd_sc_hs__a21oi_1 _5402_ (.A1(_0595_),
    .A2(_0622_),
    .B1(_0627_),
    .Y(_3587_));
 sky130_fd_sc_hs__xnor2_2 _5403_ (.A(net68),
    .B(_0598_),
    .Y(_0628_));
 sky130_fd_sc_hs__clkbuf_8 _5404_ (.A(_0107_),
    .X(_0629_));
 sky130_fd_sc_hs__nor2_1 _5405_ (.A(net108),
    .B(_0603_),
    .Y(_0630_));
 sky130_fd_sc_hs__o22ai_4 _5406_ (.A1(_0605_),
    .A2(_0573_),
    .B1(net147),
    .B2(_0427_),
    .Y(_0631_));
 sky130_fd_sc_hs__nor3_2 _5407_ (.A(_0602_),
    .B(_0630_),
    .C(_0631_),
    .Y(_0632_));
 sky130_fd_sc_hs__a21oi_4 _5408_ (.A1(net179),
    .A2(_0601_),
    .B1(_0632_),
    .Y(_0633_));
 sky130_fd_sc_hs__nor2_4 _5409_ (.A(_0629_),
    .B(_0633_),
    .Y(_0634_));
 sky130_fd_sc_hs__a21oi_2 _5410_ (.A1(_0595_),
    .A2(_0628_),
    .B1(_0634_),
    .Y(_3591_));
 sky130_fd_sc_hs__xnor2_4 _5411_ (.A(net69),
    .B(_0598_),
    .Y(_0635_));
 sky130_fd_sc_hs__nor2_1 _5412_ (.A(net110),
    .B(_0603_),
    .Y(_0636_));
 sky130_fd_sc_hs__o22ai_4 _5413_ (.A1(_0605_),
    .A2(_0574_),
    .B1(net148),
    .B2(_0427_),
    .Y(_0637_));
 sky130_fd_sc_hs__nor3_2 _5414_ (.A(_0602_),
    .B(_0636_),
    .C(_0637_),
    .Y(_0638_));
 sky130_fd_sc_hs__a21oi_4 _5415_ (.A1(net180),
    .A2(_0601_),
    .B1(_0638_),
    .Y(_0639_));
 sky130_fd_sc_hs__nor2_4 _5416_ (.A(_0629_),
    .B(_0639_),
    .Y(_0640_));
 sky130_fd_sc_hs__a21oi_2 _5417_ (.A1(_0595_),
    .A2(_0635_),
    .B1(_0640_),
    .Y(_3595_));
 sky130_fd_sc_hs__xnor2_4 _5418_ (.A(net70),
    .B(_0598_),
    .Y(_0641_));
 sky130_fd_sc_hs__nor2_1 _5419_ (.A(net116),
    .B(_0603_),
    .Y(_0642_));
 sky130_fd_sc_hs__o22ai_4 _5420_ (.A1(_0605_),
    .A2(_0575_),
    .B1(net149),
    .B2(_0427_),
    .Y(_0643_));
 sky130_fd_sc_hs__nor3_1 _5421_ (.A(_0602_),
    .B(_0642_),
    .C(_0643_),
    .Y(_0644_));
 sky130_fd_sc_hs__a21oi_2 _5422_ (.A1(net181),
    .A2(_0601_),
    .B1(_0644_),
    .Y(_0645_));
 sky130_fd_sc_hs__nor2_4 _5423_ (.A(_0629_),
    .B(_0645_),
    .Y(_0646_));
 sky130_fd_sc_hs__a21oi_2 _5424_ (.A1(_0595_),
    .A2(_0641_),
    .B1(_0646_),
    .Y(_3599_));
 sky130_fd_sc_hs__xnor2_4 _5425_ (.A(net71),
    .B(_0598_),
    .Y(_0647_));
 sky130_fd_sc_hs__nor2_1 _5426_ (.A(net117),
    .B(_0603_),
    .Y(_0648_));
 sky130_fd_sc_hs__o22ai_4 _5427_ (.A1(_0605_),
    .A2(_0576_),
    .B1(net150),
    .B2(_0427_),
    .Y(_0649_));
 sky130_fd_sc_hs__nor3_1 _5428_ (.A(_0602_),
    .B(_0648_),
    .C(_0649_),
    .Y(_0650_));
 sky130_fd_sc_hs__a21oi_1 _5429_ (.A1(net182),
    .A2(_0601_),
    .B1(_0650_),
    .Y(_0651_));
 sky130_fd_sc_hs__nor2_1 _5430_ (.A(_0629_),
    .B(_0651_),
    .Y(_0652_));
 sky130_fd_sc_hs__a21oi_2 _5431_ (.A1(_0595_),
    .A2(_0647_),
    .B1(_0652_),
    .Y(_3603_));
 sky130_fd_sc_hs__clkbuf_8 _5432_ (.A(_0108_),
    .X(_0653_));
 sky130_fd_sc_hs__xnor2_4 _5433_ (.A(net72),
    .B(_0598_),
    .Y(_0654_));
 sky130_fd_sc_hs__nor2_1 _5434_ (.A(net118),
    .B(_0603_),
    .Y(_0655_));
 sky130_fd_sc_hs__o22ai_4 _5435_ (.A1(_0605_),
    .A2(_0577_),
    .B1(net151),
    .B2(_0427_),
    .Y(_0656_));
 sky130_fd_sc_hs__nor3_1 _5436_ (.A(_0602_),
    .B(_0655_),
    .C(_0656_),
    .Y(_0657_));
 sky130_fd_sc_hs__a21oi_2 _5437_ (.A1(net183),
    .A2(_0601_),
    .B1(_0657_),
    .Y(_0658_));
 sky130_fd_sc_hs__nor2_1 _5438_ (.A(_0629_),
    .B(_0658_),
    .Y(_0659_));
 sky130_fd_sc_hs__a21oi_2 _5439_ (.A1(_0653_),
    .A2(_0654_),
    .B1(_0659_),
    .Y(_3607_));
 sky130_fd_sc_hs__xnor2_4 _5440_ (.A(net73),
    .B(_0598_),
    .Y(_0660_));
 sky130_fd_sc_hs__buf_4 _5441_ (.A(net366),
    .X(_0661_));
 sky130_fd_sc_hs__nor2_1 _5442_ (.A(net119),
    .B(_0603_),
    .Y(_0662_));
 sky130_fd_sc_hs__buf_8 _5443_ (.A(_0383_),
    .X(_0663_));
 sky130_fd_sc_hs__o22ai_4 _5444_ (.A1(_0605_),
    .A2(_0578_),
    .B1(net152),
    .B2(_0663_),
    .Y(_0664_));
 sky130_fd_sc_hs__nor3_1 _5445_ (.A(_0661_),
    .B(_0662_),
    .C(_0664_),
    .Y(_0665_));
 sky130_fd_sc_hs__a21oi_2 _5446_ (.A1(net184),
    .A2(_0601_),
    .B1(_0665_),
    .Y(_0666_));
 sky130_fd_sc_hs__nor2_4 _5447_ (.A(_0629_),
    .B(_0666_),
    .Y(_0667_));
 sky130_fd_sc_hs__a21oi_1 _5448_ (.A1(_0653_),
    .A2(_0660_),
    .B1(_0667_),
    .Y(_3611_));
 sky130_fd_sc_hs__buf_16 _5449_ (.A(_0597_),
    .X(_0668_));
 sky130_fd_sc_hs__xnor2_2 _5450_ (.A(net43),
    .B(_0668_),
    .Y(_0669_));
 sky130_fd_sc_hs__clkbuf_8 _5451_ (.A(_0379_),
    .X(_0670_));
 sky130_fd_sc_hs__clkbuf_4 _5452_ (.A(_0387_),
    .X(_0671_));
 sky130_fd_sc_hs__nor2_1 _5453_ (.A(net82),
    .B(_0671_),
    .Y(_0672_));
 sky130_fd_sc_hs__buf_8 _5454_ (.A(_0381_),
    .X(_0673_));
 sky130_fd_sc_hs__o22ai_4 _5455_ (.A1(_0673_),
    .A2(_0580_),
    .B1(net122),
    .B2(_0663_),
    .Y(_0674_));
 sky130_fd_sc_hs__nor3_1 _5456_ (.A(_0661_),
    .B(_0672_),
    .C(_0674_),
    .Y(_0675_));
 sky130_fd_sc_hs__a21oi_2 _5457_ (.A1(net154),
    .A2(_0670_),
    .B1(_0675_),
    .Y(_0676_));
 sky130_fd_sc_hs__nor2_2 _5458_ (.A(_0629_),
    .B(_0676_),
    .Y(_0677_));
 sky130_fd_sc_hs__a21oi_1 _5459_ (.A1(_0653_),
    .A2(_0669_),
    .B1(_0677_),
    .Y(_3615_));
 sky130_fd_sc_hs__xnor2_4 _5460_ (.A(net44),
    .B(_0668_),
    .Y(_0678_));
 sky130_fd_sc_hs__nor2_1 _5461_ (.A(net83),
    .B(_0671_),
    .Y(_0679_));
 sky130_fd_sc_hs__o22ai_2 _5462_ (.A1(_0673_),
    .A2(_0581_),
    .B1(net123),
    .B2(_0663_),
    .Y(_0680_));
 sky130_fd_sc_hs__nor3_2 _5463_ (.A(_0661_),
    .B(_0679_),
    .C(_0680_),
    .Y(_0681_));
 sky130_fd_sc_hs__a21oi_4 _5464_ (.A1(net155),
    .A2(_0670_),
    .B1(_0681_),
    .Y(_0682_));
 sky130_fd_sc_hs__nor2_2 _5465_ (.A(_0629_),
    .B(_0682_),
    .Y(_0683_));
 sky130_fd_sc_hs__a21oi_1 _5466_ (.A1(_0653_),
    .A2(_0678_),
    .B1(_0683_),
    .Y(_3619_));
 sky130_fd_sc_hs__xnor2_4 _5467_ (.A(net45),
    .B(_0668_),
    .Y(_0684_));
 sky130_fd_sc_hs__nor2_1 _5468_ (.A(net84),
    .B(_0671_),
    .Y(_0685_));
 sky130_fd_sc_hs__o22ai_1 _5469_ (.A1(_0673_),
    .A2(_0582_),
    .B1(net124),
    .B2(_0663_),
    .Y(_0686_));
 sky130_fd_sc_hs__nor3_1 _5470_ (.A(_0661_),
    .B(_0685_),
    .C(_0686_),
    .Y(_0687_));
 sky130_fd_sc_hs__a21oi_2 _5471_ (.A1(net156),
    .A2(_0670_),
    .B1(_0687_),
    .Y(_0688_));
 sky130_fd_sc_hs__nor2_1 _5472_ (.A(_0629_),
    .B(_0688_),
    .Y(_0689_));
 sky130_fd_sc_hs__a21oi_2 _5473_ (.A1(_0653_),
    .A2(_0684_),
    .B1(_0689_),
    .Y(_3623_));
 sky130_fd_sc_hs__xnor2_4 _5474_ (.A(net46),
    .B(_0668_),
    .Y(_0690_));
 sky130_fd_sc_hs__nor2_1 _5475_ (.A(net85),
    .B(_0671_),
    .Y(_0691_));
 sky130_fd_sc_hs__o22ai_2 _5476_ (.A1(_0673_),
    .A2(_0584_),
    .B1(net125),
    .B2(_0663_),
    .Y(_0692_));
 sky130_fd_sc_hs__nor3_1 _5477_ (.A(_0661_),
    .B(_0691_),
    .C(_0692_),
    .Y(_0693_));
 sky130_fd_sc_hs__a21oi_2 _5478_ (.A1(net157),
    .A2(_0670_),
    .B1(_0693_),
    .Y(_0694_));
 sky130_fd_sc_hs__nor2_1 _5479_ (.A(_0629_),
    .B(_0694_),
    .Y(_0695_));
 sky130_fd_sc_hs__a21oi_2 _5480_ (.A1(_0653_),
    .A2(_0690_),
    .B1(_0695_),
    .Y(_3627_));
 sky130_fd_sc_hs__xnor2_4 _5481_ (.A(net47),
    .B(_0668_),
    .Y(_0696_));
 sky130_fd_sc_hs__buf_4 _5482_ (.A(_0107_),
    .X(_0697_));
 sky130_fd_sc_hs__nor2_1 _5483_ (.A(net86),
    .B(_0671_),
    .Y(_0698_));
 sky130_fd_sc_hs__o22ai_2 _5484_ (.A1(_0673_),
    .A2(_0585_),
    .B1(net126),
    .B2(_0663_),
    .Y(_0699_));
 sky130_fd_sc_hs__nor3_1 _5485_ (.A(_0661_),
    .B(_0698_),
    .C(_0699_),
    .Y(_0700_));
 sky130_fd_sc_hs__a21oi_2 _5486_ (.A1(net158),
    .A2(_0670_),
    .B1(_0700_),
    .Y(_0701_));
 sky130_fd_sc_hs__nor2_1 _5487_ (.A(_0697_),
    .B(_0701_),
    .Y(_0702_));
 sky130_fd_sc_hs__a21oi_1 _5488_ (.A1(_0653_),
    .A2(_0696_),
    .B1(_0702_),
    .Y(_3631_));
 sky130_fd_sc_hs__xnor2_4 _5489_ (.A(net48),
    .B(_0668_),
    .Y(_0703_));
 sky130_fd_sc_hs__nor2_1 _5490_ (.A(net87),
    .B(_0671_),
    .Y(_0704_));
 sky130_fd_sc_hs__o22ai_2 _5491_ (.A1(_0673_),
    .A2(net107),
    .B1(net127),
    .B2(_0663_),
    .Y(_0705_));
 sky130_fd_sc_hs__nor3_1 _5492_ (.A(_0661_),
    .B(_0704_),
    .C(_0705_),
    .Y(_0706_));
 sky130_fd_sc_hs__a21oi_1 _5493_ (.A1(net159),
    .A2(_0670_),
    .B1(_0706_),
    .Y(_0707_));
 sky130_fd_sc_hs__nor2_1 _5494_ (.A(_0697_),
    .B(_0707_),
    .Y(_0708_));
 sky130_fd_sc_hs__a21oi_1 _5495_ (.A1(_0653_),
    .A2(_0703_),
    .B1(_0708_),
    .Y(_3635_));
 sky130_fd_sc_hs__xnor2_4 _5496_ (.A(net49),
    .B(_0668_),
    .Y(_0709_));
 sky130_fd_sc_hs__nor2_1 _5497_ (.A(net88),
    .B(_0671_),
    .Y(_0710_));
 sky130_fd_sc_hs__o22ai_2 _5498_ (.A1(_0673_),
    .A2(_0436_),
    .B1(net128),
    .B2(_0663_),
    .Y(_0711_));
 sky130_fd_sc_hs__nor3_1 _5499_ (.A(_0661_),
    .B(_0710_),
    .C(_0711_),
    .Y(_0712_));
 sky130_fd_sc_hs__a21oi_1 _5500_ (.A1(net160),
    .A2(_0670_),
    .B1(_0712_),
    .Y(_0713_));
 sky130_fd_sc_hs__nor2_1 _5501_ (.A(_0697_),
    .B(_0713_),
    .Y(_0714_));
 sky130_fd_sc_hs__a21oi_1 _5502_ (.A1(_0653_),
    .A2(_0709_),
    .B1(_0714_),
    .Y(_3639_));
 sky130_fd_sc_hs__xnor2_4 _5503_ (.A(net50),
    .B(_0668_),
    .Y(_0715_));
 sky130_fd_sc_hs__nor2_1 _5504_ (.A(net89),
    .B(_0671_),
    .Y(_0716_));
 sky130_fd_sc_hs__o22ai_2 _5505_ (.A1(_0673_),
    .A2(_0446_),
    .B1(net129),
    .B2(_0663_),
    .Y(_0717_));
 sky130_fd_sc_hs__nor3_1 _5506_ (.A(_0661_),
    .B(_0716_),
    .C(_0717_),
    .Y(_0718_));
 sky130_fd_sc_hs__a21oi_1 _5507_ (.A1(net161),
    .A2(_0670_),
    .B1(_0718_),
    .Y(_0719_));
 sky130_fd_sc_hs__nor2_1 _5508_ (.A(_0697_),
    .B(_0719_),
    .Y(_0720_));
 sky130_fd_sc_hs__a21oi_1 _5509_ (.A1(_0653_),
    .A2(_0715_),
    .B1(_0720_),
    .Y(_3643_));
 sky130_fd_sc_hs__buf_4 _5510_ (.A(_0107_),
    .X(_0721_));
 sky130_fd_sc_hs__xnor2_4 _5511_ (.A(net51),
    .B(_0668_),
    .Y(_0722_));
 sky130_fd_sc_hs__nor2_1 _5512_ (.A(net90),
    .B(_0671_),
    .Y(_0723_));
 sky130_fd_sc_hs__o22ai_2 _5513_ (.A1(_0673_),
    .A2(_0449_),
    .B1(net130),
    .B2(_0663_),
    .Y(_0724_));
 sky130_fd_sc_hs__nor3_1 _5514_ (.A(_0661_),
    .B(_0723_),
    .C(_0724_),
    .Y(_0725_));
 sky130_fd_sc_hs__a21oi_1 _5515_ (.A1(net162),
    .A2(_0670_),
    .B1(_0725_),
    .Y(_0726_));
 sky130_fd_sc_hs__nor2_1 _5516_ (.A(_0697_),
    .B(_0726_),
    .Y(_0727_));
 sky130_fd_sc_hs__a21oi_1 _5517_ (.A1(_0721_),
    .A2(_0722_),
    .B1(_0727_),
    .Y(_3647_));
 sky130_fd_sc_hs__xnor2_4 _5518_ (.A(net52),
    .B(_0668_),
    .Y(_0728_));
 sky130_fd_sc_hs__clkbuf_8 _5519_ (.A(net366),
    .X(_0729_));
 sky130_fd_sc_hs__nor2_1 _5520_ (.A(net91),
    .B(_0671_),
    .Y(_0730_));
 sky130_fd_sc_hs__buf_8 _5521_ (.A(_0383_),
    .X(_0731_));
 sky130_fd_sc_hs__o22ai_4 _5522_ (.A1(_0673_),
    .A2(_0586_),
    .B1(net131),
    .B2(_0731_),
    .Y(_0732_));
 sky130_fd_sc_hs__nor3_1 _5523_ (.A(_0729_),
    .B(_0730_),
    .C(_0732_),
    .Y(_0733_));
 sky130_fd_sc_hs__a21oi_1 _5524_ (.A1(net163),
    .A2(_0670_),
    .B1(_0733_),
    .Y(_0734_));
 sky130_fd_sc_hs__nor2_2 _5525_ (.A(_0697_),
    .B(_0734_),
    .Y(_0735_));
 sky130_fd_sc_hs__a21oi_1 _5526_ (.A1(_0721_),
    .A2(_0728_),
    .B1(_0735_),
    .Y(_3651_));
 sky130_fd_sc_hs__buf_8 _5527_ (.A(_0597_),
    .X(_0736_));
 sky130_fd_sc_hs__xnor2_4 _5528_ (.A(net54),
    .B(_0736_),
    .Y(_0737_));
 sky130_fd_sc_hs__clkbuf_16 _5529_ (.A(net366),
    .X(_0738_));
 sky130_fd_sc_hs__buf_4 _5530_ (.A(_0387_),
    .X(_0739_));
 sky130_fd_sc_hs__nor2_1 _5531_ (.A(net93),
    .B(_0739_),
    .Y(_0740_));
 sky130_fd_sc_hs__buf_8 _5532_ (.A(_0381_),
    .X(_0741_));
 sky130_fd_sc_hs__o22ai_4 _5533_ (.A1(_0741_),
    .A2(_0588_),
    .B1(net133),
    .B2(_0731_),
    .Y(_0742_));
 sky130_fd_sc_hs__nor3_2 _5534_ (.A(_0729_),
    .B(_0740_),
    .C(_0742_),
    .Y(_0743_));
 sky130_fd_sc_hs__a21oi_4 _5535_ (.A1(net165),
    .A2(_0738_),
    .B1(_0743_),
    .Y(_0744_));
 sky130_fd_sc_hs__nor2_2 _5536_ (.A(_0697_),
    .B(_0744_),
    .Y(_0745_));
 sky130_fd_sc_hs__a21oi_1 _5537_ (.A1(_0721_),
    .A2(_0737_),
    .B1(_0745_),
    .Y(_3655_));
 sky130_fd_sc_hs__xnor2_2 _5538_ (.A(net55),
    .B(_0736_),
    .Y(_0746_));
 sky130_fd_sc_hs__nor2_1 _5539_ (.A(net94),
    .B(_0739_),
    .Y(_0747_));
 sky130_fd_sc_hs__o22ai_4 _5540_ (.A1(_0741_),
    .A2(net109),
    .B1(net134),
    .B2(_0731_),
    .Y(_0748_));
 sky130_fd_sc_hs__nor3_2 _5541_ (.A(_0729_),
    .B(_0747_),
    .C(_0748_),
    .Y(_0749_));
 sky130_fd_sc_hs__a21oi_4 _5542_ (.A1(net166),
    .A2(_0738_),
    .B1(_0749_),
    .Y(_0750_));
 sky130_fd_sc_hs__nor2_2 _5543_ (.A(_0697_),
    .B(_0750_),
    .Y(_0751_));
 sky130_fd_sc_hs__a21oi_1 _5544_ (.A1(_0721_),
    .A2(_0746_),
    .B1(_0751_),
    .Y(_3659_));
 sky130_fd_sc_hs__xnor2_1 _5545_ (.A(net56),
    .B(_0736_),
    .Y(_0752_));
 sky130_fd_sc_hs__nor2_1 _5546_ (.A(net95),
    .B(_0739_),
    .Y(_0753_));
 sky130_fd_sc_hs__o22ai_4 _5547_ (.A1(_0741_),
    .A2(_0520_),
    .B1(net135),
    .B2(_0731_),
    .Y(_0754_));
 sky130_fd_sc_hs__nor3_2 _5548_ (.A(_0729_),
    .B(_0753_),
    .C(_0754_),
    .Y(_0755_));
 sky130_fd_sc_hs__a21oi_4 _5549_ (.A1(net167),
    .A2(_0738_),
    .B1(_0755_),
    .Y(_0756_));
 sky130_fd_sc_hs__nor2_4 _5550_ (.A(_0697_),
    .B(_0756_),
    .Y(_0757_));
 sky130_fd_sc_hs__a21oi_1 _5551_ (.A1(_0721_),
    .A2(_0752_),
    .B1(_0757_),
    .Y(_3663_));
 sky130_fd_sc_hs__xnor2_1 _5552_ (.A(net57),
    .B(_0736_),
    .Y(_0758_));
 sky130_fd_sc_hs__nor2_1 _5553_ (.A(net96),
    .B(_0739_),
    .Y(_0759_));
 sky130_fd_sc_hs__o22ai_4 _5554_ (.A1(_0741_),
    .A2(_0526_),
    .B1(net136),
    .B2(_0731_),
    .Y(_0760_));
 sky130_fd_sc_hs__nor3_2 _5555_ (.A(_0729_),
    .B(_0759_),
    .C(_0760_),
    .Y(_0761_));
 sky130_fd_sc_hs__a21oi_4 _5556_ (.A1(net168),
    .A2(_0738_),
    .B1(_0761_),
    .Y(_0762_));
 sky130_fd_sc_hs__nor2_4 _5557_ (.A(_0697_),
    .B(_0762_),
    .Y(_0763_));
 sky130_fd_sc_hs__a21oi_1 _5558_ (.A1(_0721_),
    .A2(_0758_),
    .B1(_0763_),
    .Y(_3667_));
 sky130_fd_sc_hs__xnor2_1 _5559_ (.A(net58),
    .B(_0736_),
    .Y(_0764_));
 sky130_fd_sc_hs__nor2_1 _5560_ (.A(net97),
    .B(_0739_),
    .Y(_0765_));
 sky130_fd_sc_hs__o22ai_4 _5561_ (.A1(_0741_),
    .A2(_0527_),
    .B1(net137),
    .B2(_0731_),
    .Y(_0766_));
 sky130_fd_sc_hs__nor3_2 _5562_ (.A(_0729_),
    .B(_0765_),
    .C(_0766_),
    .Y(_0767_));
 sky130_fd_sc_hs__a21oi_4 _5563_ (.A1(net169),
    .A2(_0738_),
    .B1(_0767_),
    .Y(_0768_));
 sky130_fd_sc_hs__nor2_1 _5564_ (.A(_0568_),
    .B(_0768_),
    .Y(_0769_));
 sky130_fd_sc_hs__a21oi_2 _5565_ (.A1(_0721_),
    .A2(_0764_),
    .B1(_0769_),
    .Y(_3671_));
 sky130_fd_sc_hs__xnor2_2 _5566_ (.A(net59),
    .B(_0736_),
    .Y(_0770_));
 sky130_fd_sc_hs__nor2_1 _5567_ (.A(net98),
    .B(_0739_),
    .Y(_0771_));
 sky130_fd_sc_hs__o22ai_4 _5568_ (.A1(_0741_),
    .A2(_0529_),
    .B1(net138),
    .B2(_0731_),
    .Y(_0772_));
 sky130_fd_sc_hs__nor3_2 _5569_ (.A(_0729_),
    .B(_0771_),
    .C(_0772_),
    .Y(_0773_));
 sky130_fd_sc_hs__a21oi_4 _5570_ (.A1(net170),
    .A2(_0738_),
    .B1(_0773_),
    .Y(_0774_));
 sky130_fd_sc_hs__nor2_1 _5571_ (.A(_0568_),
    .B(_0774_),
    .Y(_0775_));
 sky130_fd_sc_hs__a21oi_2 _5572_ (.A1(_0721_),
    .A2(_0770_),
    .B1(_0775_),
    .Y(_3675_));
 sky130_fd_sc_hs__xnor2_1 _5573_ (.A(net60),
    .B(_0736_),
    .Y(_0776_));
 sky130_fd_sc_hs__nor2_1 _5574_ (.A(net99),
    .B(_0739_),
    .Y(_0777_));
 sky130_fd_sc_hs__o22ai_4 _5575_ (.A1(_0741_),
    .A2(_0565_),
    .B1(net139),
    .B2(_0731_),
    .Y(_0778_));
 sky130_fd_sc_hs__nor3_2 _5576_ (.A(_0729_),
    .B(_0777_),
    .C(_0778_),
    .Y(_0779_));
 sky130_fd_sc_hs__a21oi_4 _5577_ (.A1(net171),
    .A2(_0738_),
    .B1(_0779_),
    .Y(_0780_));
 sky130_fd_sc_hs__nor2_1 _5578_ (.A(_0568_),
    .B(_0780_),
    .Y(_0781_));
 sky130_fd_sc_hs__a21oi_1 _5579_ (.A1(_0721_),
    .A2(_0776_),
    .B1(_0781_),
    .Y(_3679_));
 sky130_fd_sc_hs__xnor2_1 _5580_ (.A(net61),
    .B(_0736_),
    .Y(_0782_));
 sky130_fd_sc_hs__nor2_1 _5581_ (.A(net100),
    .B(_0739_),
    .Y(_0783_));
 sky130_fd_sc_hs__o22ai_2 _5582_ (.A1(_0741_),
    .A2(_0566_),
    .B1(net140),
    .B2(_0731_),
    .Y(_0784_));
 sky130_fd_sc_hs__nor3_2 _5583_ (.A(_0729_),
    .B(_0783_),
    .C(_0784_),
    .Y(_0785_));
 sky130_fd_sc_hs__a21oi_4 _5584_ (.A1(net172),
    .A2(_0738_),
    .B1(_0785_),
    .Y(_0786_));
 sky130_fd_sc_hs__nor2_1 _5585_ (.A(_0568_),
    .B(_0786_),
    .Y(_0787_));
 sky130_fd_sc_hs__a21oi_1 _5586_ (.A1(_0721_),
    .A2(_0782_),
    .B1(_0787_),
    .Y(_3683_));
 sky130_fd_sc_hs__buf_8 _5587_ (.A(_0107_),
    .X(_0788_));
 sky130_fd_sc_hs__xnor2_1 _5588_ (.A(net62),
    .B(_0736_),
    .Y(_0789_));
 sky130_fd_sc_hs__nor2_1 _5589_ (.A(net101),
    .B(_0739_),
    .Y(_0790_));
 sky130_fd_sc_hs__o22ai_2 _5590_ (.A1(_0741_),
    .A2(net111),
    .B1(net141),
    .B2(_0731_),
    .Y(_0791_));
 sky130_fd_sc_hs__nor3_2 _5591_ (.A(_0729_),
    .B(_0790_),
    .C(_0791_),
    .Y(_0792_));
 sky130_fd_sc_hs__a21oi_4 _5592_ (.A1(net173),
    .A2(_0738_),
    .B1(_0792_),
    .Y(_0793_));
 sky130_fd_sc_hs__nor2_1 _5593_ (.A(_0568_),
    .B(_0793_),
    .Y(_0794_));
 sky130_fd_sc_hs__a21oi_1 _5594_ (.A1(_0788_),
    .A2(_0789_),
    .B1(_0794_),
    .Y(_3687_));
 sky130_fd_sc_hs__xnor2_1 _5595_ (.A(net63),
    .B(_0736_),
    .Y(_0795_));
 sky130_fd_sc_hs__nor2_1 _5596_ (.A(net102),
    .B(_0739_),
    .Y(_0796_));
 sky130_fd_sc_hs__o22ai_4 _5597_ (.A1(_0741_),
    .A2(net112),
    .B1(net142),
    .B2(_0383_),
    .Y(_0797_));
 sky130_fd_sc_hs__nor3_2 _5598_ (.A(net366),
    .B(_0796_),
    .C(_0797_),
    .Y(_0798_));
 sky130_fd_sc_hs__a21oi_4 _5599_ (.A1(net174),
    .A2(_0738_),
    .B1(_0798_),
    .Y(_0799_));
 sky130_fd_sc_hs__nor2_1 _5600_ (.A(_0568_),
    .B(_0799_),
    .Y(_0800_));
 sky130_fd_sc_hs__a21oi_1 _5601_ (.A1(_0788_),
    .A2(_0795_),
    .B1(_0800_),
    .Y(_3691_));
 sky130_fd_sc_hs__xnor2_2 _5602_ (.A(net65),
    .B(_0597_),
    .Y(_0801_));
 sky130_fd_sc_hs__nor2_1 _5603_ (.A(net104),
    .B(_0387_),
    .Y(_0802_));
 sky130_fd_sc_hs__o22ai_4 _5604_ (.A1(_0381_),
    .A2(_0567_),
    .B1(net144),
    .B2(_0383_),
    .Y(_0803_));
 sky130_fd_sc_hs__nor3_2 _5605_ (.A(net366),
    .B(_0802_),
    .C(_0803_),
    .Y(_0804_));
 sky130_fd_sc_hs__a21oi_4 _5606_ (.A1(net176),
    .A2(_0602_),
    .B1(_0804_),
    .Y(_0805_));
 sky130_fd_sc_hs__nor2_1 _5607_ (.A(_0568_),
    .B(_0805_),
    .Y(_0806_));
 sky130_fd_sc_hs__a21oi_1 _5608_ (.A1(_0788_),
    .A2(_0801_),
    .B1(_0806_),
    .Y(_3695_));
 sky130_fd_sc_hs__inv_2 _5609_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .Y(_3703_));
 sky130_fd_sc_hs__inv_1 _5610_ (.A(_2234_),
    .Y(_3714_));
 sky130_fd_sc_hs__inv_1 _5611_ (.A(_2239_),
    .Y(_2242_));
 sky130_fd_sc_hs__nand2b_4 _5612_ (.A_N(\genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[2] ),
    .B(_0087_),
    .Y(_0807_));
 sky130_fd_sc_hs__clkbuf_4 _5613_ (.A(_0807_),
    .X(_0808_));
 sky130_fd_sc_hs__a22o_1 _5614_ (.A1(_0572_),
    .A2(_0086_),
    .B1(_0808_),
    .B2(_0586_),
    .X(_2247_));
 sky130_fd_sc_hs__inv_1 _5615_ (.A(_2253_),
    .Y(_3722_));
 sky130_fd_sc_hs__a22o_1 _5616_ (.A1(_0573_),
    .A2(_0086_),
    .B1(_0808_),
    .B2(_0588_),
    .X(_2256_));
 sky130_fd_sc_hs__inv_1 _5617_ (.A(_2268_),
    .Y(_2271_));
 sky130_fd_sc_hs__clkbuf_4 _5618_ (.A(_0085_),
    .X(_0809_));
 sky130_fd_sc_hs__a22o_1 _5619_ (.A1(_0574_),
    .A2(_0809_),
    .B1(_0808_),
    .B2(net109),
    .X(_2276_));
 sky130_fd_sc_hs__inv_1 _5620_ (.A(_2290_),
    .Y(_3733_));
 sky130_fd_sc_hs__a22o_1 _5621_ (.A1(_0575_),
    .A2(_0809_),
    .B1(_0808_),
    .B2(_0520_),
    .X(_2293_));
 sky130_fd_sc_hs__inv_1 _5622_ (.A(_2311_),
    .Y(_3745_));
 sky130_fd_sc_hs__a22o_1 _5623_ (.A1(_0576_),
    .A2(_0809_),
    .B1(_0808_),
    .B2(_0526_),
    .X(_2315_));
 sky130_fd_sc_hs__inv_1 _5624_ (.A(_2341_),
    .Y(_3751_));
 sky130_fd_sc_hs__a22o_1 _5625_ (.A1(_0577_),
    .A2(_0809_),
    .B1(_0808_),
    .B2(_0527_),
    .X(_2350_));
 sky130_fd_sc_hs__inv_1 _5626_ (.A(_2375_),
    .Y(_3760_));
 sky130_fd_sc_hs__a22o_2 _5627_ (.A1(_0578_),
    .A2(_0809_),
    .B1(_0808_),
    .B2(_0529_),
    .X(_2378_));
 sky130_fd_sc_hs__inv_1 _5628_ (.A(_2406_),
    .Y(_3773_));
 sky130_fd_sc_hs__a22o_2 _5629_ (.A1(_0580_),
    .A2(_0809_),
    .B1(_0808_),
    .B2(_0565_),
    .X(_2410_));
 sky130_fd_sc_hs__a22o_2 _5630_ (.A1(_0581_),
    .A2(_0809_),
    .B1(_0808_),
    .B2(_0566_),
    .X(_2448_));
 sky130_fd_sc_hs__inv_1 _5631_ (.A(_2431_),
    .Y(_2482_));
 sky130_fd_sc_hs__a22o_2 _5632_ (.A1(_0582_),
    .A2(_0809_),
    .B1(_0808_),
    .B2(net111),
    .X(_2493_));
 sky130_fd_sc_hs__inv_1 _5633_ (.A(_2532_),
    .Y(_2534_));
 sky130_fd_sc_hs__a22o_2 _5634_ (.A1(_0584_),
    .A2(_0809_),
    .B1(_0807_),
    .B2(net112),
    .X(_2539_));
 sky130_fd_sc_hs__inv_1 _5635_ (.A(_2514_),
    .Y(_2581_));
 sky130_fd_sc_hs__inv_1 _5636_ (.A(_2586_),
    .Y(_2589_));
 sky130_fd_sc_hs__inv_1 _5637_ (.A(_2529_),
    .Y(_3802_));
 sky130_fd_sc_hs__a22o_2 _5638_ (.A1(_0585_),
    .A2(_0809_),
    .B1(_0807_),
    .B2(_0567_),
    .X(_2594_));
 sky130_fd_sc_hs__inv_1 _5639_ (.A(_2560_),
    .Y(_2636_));
 sky130_fd_sc_hs__inv_1 _5640_ (.A(_2648_),
    .Y(_3811_));
 sky130_fd_sc_hs__a22o_2 _5641_ (.A1(net107),
    .A2(_0085_),
    .B1(_0807_),
    .B2(_0382_),
    .X(_2652_));
 sky130_fd_sc_hs__inv_1 _5642_ (.A(_2701_),
    .Y(_3822_));
 sky130_fd_sc_hs__inv_1 _5643_ (.A(_2692_),
    .Y(_2764_));
 sky130_fd_sc_hs__inv_1 _5644_ (.A(_2772_),
    .Y(_3826_));
 sky130_fd_sc_hs__inv_1 _5645_ (.A(_2830_),
    .Y(_3829_));
 sky130_fd_sc_hs__inv_1 _5646_ (.A(_2838_),
    .Y(_3832_));
 sky130_fd_sc_hs__inv_1 _5647_ (.A(_2892_),
    .Y(_3836_));
 sky130_fd_sc_hs__inv_1 _5648_ (.A(_2817_),
    .Y(_2895_));
 sky130_fd_sc_hs__inv_1 _5649_ (.A(_2902_),
    .Y(_3838_));
 sky130_fd_sc_hs__inv_1 _5650_ (.A(_2955_),
    .Y(_3842_));
 sky130_fd_sc_hs__inv_1 _5651_ (.A(_2879_),
    .Y(_2958_));
 sky130_fd_sc_hs__inv_1 _5652_ (.A(_2966_),
    .Y(_3844_));
 sky130_fd_sc_hs__inv_1 _5653_ (.A(_3018_),
    .Y(_3848_));
 sky130_fd_sc_hs__inv_1 _5654_ (.A(_2942_),
    .Y(_3021_));
 sky130_fd_sc_hs__inv_1 _5655_ (.A(_3029_),
    .Y(_3850_));
 sky130_fd_sc_hs__inv_1 _5656_ (.A(_3077_),
    .Y(_3854_));
 sky130_fd_sc_hs__inv_1 _5657_ (.A(_3005_),
    .Y(_3080_));
 sky130_fd_sc_hs__inv_1 _5658_ (.A(_3088_),
    .Y(_3856_));
 sky130_fd_sc_hs__inv_1 _5659_ (.A(_3134_),
    .Y(_3860_));
 sky130_fd_sc_hs__inv_1 _5660_ (.A(_3064_),
    .Y(_3137_));
 sky130_fd_sc_hs__inv_1 _5661_ (.A(_3145_),
    .Y(_3862_));
 sky130_fd_sc_hs__inv_1 _5662_ (.A(_3192_),
    .Y(_3866_));
 sky130_fd_sc_hs__inv_1 _5663_ (.A(_3121_),
    .Y(_3195_));
 sky130_fd_sc_hs__inv_1 _5664_ (.A(_3203_),
    .Y(_3868_));
 sky130_fd_sc_hs__inv_1 _5665_ (.A(_3246_),
    .Y(_3872_));
 sky130_fd_sc_hs__inv_1 _5666_ (.A(_3179_),
    .Y(_3249_));
 sky130_fd_sc_hs__inv_1 _5667_ (.A(_3257_),
    .Y(_3874_));
 sky130_fd_sc_hs__inv_1 _5668_ (.A(_3296_),
    .Y(_3878_));
 sky130_fd_sc_hs__inv_1 _5669_ (.A(_3233_),
    .Y(_3299_));
 sky130_fd_sc_hs__inv_1 _5670_ (.A(_3307_),
    .Y(_3880_));
 sky130_fd_sc_hs__inv_1 _5671_ (.A(_3310_),
    .Y(_3311_));
 sky130_fd_sc_hs__inv_1 _5672_ (.A(_3345_),
    .Y(_3884_));
 sky130_fd_sc_hs__inv_1 _5673_ (.A(_3282_),
    .Y(_3348_));
 sky130_fd_sc_hs__inv_1 _5674_ (.A(_3356_),
    .Y(_3886_));
 sky130_fd_sc_hs__inv_1 _5675_ (.A(_3388_),
    .Y(_3890_));
 sky130_fd_sc_hs__inv_1 _5676_ (.A(_3330_),
    .Y(_3391_));
 sky130_fd_sc_hs__inv_1 _5677_ (.A(_3399_),
    .Y(_3892_));
 sky130_fd_sc_hs__inv_1 _5678_ (.A(_3213_),
    .Y(_3265_));
 sky130_fd_sc_hs__inv_1 _5679_ (.A(_3427_),
    .Y(_3896_));
 sky130_fd_sc_hs__inv_1 _5680_ (.A(_3438_),
    .Y(_3898_));
 sky130_fd_sc_hs__inv_1 _5681_ (.A(_3465_),
    .Y(_3902_));
 sky130_fd_sc_hs__inv_1 _5682_ (.A(_3414_),
    .Y(_3468_));
 sky130_fd_sc_hs__inv_1 _5683_ (.A(_3476_),
    .Y(_3904_));
 sky130_fd_sc_hs__inv_1 _5684_ (.A(_3483_),
    .Y(_3488_));
 sky130_fd_sc_hs__inv_1 _5685_ (.A(_3500_),
    .Y(_3908_));
 sky130_fd_sc_hs__inv_1 _5686_ (.A(_3452_),
    .Y(_3503_));
 sky130_fd_sc_hs__inv_1 _5687_ (.A(_3512_),
    .Y(_3910_));
 sky130_fd_sc_hs__inv_1 _5688_ (.A(_3529_),
    .Y(_3914_));
 sky130_fd_sc_hs__inv_1 _5689_ (.A(_3541_),
    .Y(_3916_));
 sky130_fd_sc_hs__inv_1 _5690_ (.A(_3484_),
    .Y(_3532_));
 sky130_fd_sc_hs__inv_1 _5691_ (.A(_3565_),
    .Y(_3924_));
 sky130_fd_sc_hs__inv_1 _5692_ (.A(net66),
    .Y(_3928_));
 sky130_fd_sc_hs__inv_1 _5693_ (.A(net69),
    .Y(_3966_));
 sky130_fd_sc_hs__inv_1 _5694_ (.A(net70),
    .Y(_3972_));
 sky130_fd_sc_hs__inv_1 _5695_ (.A(net71),
    .Y(_3978_));
 sky130_fd_sc_hs__inv_1 _5696_ (.A(net72),
    .Y(_3984_));
 sky130_fd_sc_hs__inv_1 _5697_ (.A(net73),
    .Y(_3990_));
 sky130_fd_sc_hs__inv_1 _5698_ (.A(net43),
    .Y(_3996_));
 sky130_fd_sc_hs__inv_1 _5699_ (.A(net44),
    .Y(_4002_));
 sky130_fd_sc_hs__inv_1 _5700_ (.A(net45),
    .Y(_4008_));
 sky130_fd_sc_hs__inv_1 _5701_ (.A(net46),
    .Y(_4014_));
 sky130_fd_sc_hs__inv_1 _5702_ (.A(net47),
    .Y(_4020_));
 sky130_fd_sc_hs__inv_1 _5703_ (.A(net48),
    .Y(_4026_));
 sky130_fd_sc_hs__inv_1 _5704_ (.A(net49),
    .Y(_4032_));
 sky130_fd_sc_hs__inv_1 _5705_ (.A(net50),
    .Y(_4038_));
 sky130_fd_sc_hs__inv_1 _5706_ (.A(net51),
    .Y(_4044_));
 sky130_fd_sc_hs__inv_1 _5707_ (.A(net52),
    .Y(_4050_));
 sky130_fd_sc_hs__inv_1 _5708_ (.A(net54),
    .Y(_4056_));
 sky130_fd_sc_hs__inv_1 _5709_ (.A(net55),
    .Y(_4062_));
 sky130_fd_sc_hs__inv_1 _5710_ (.A(net56),
    .Y(_4068_));
 sky130_fd_sc_hs__inv_1 _5711_ (.A(net57),
    .Y(_4074_));
 sky130_fd_sc_hs__inv_1 _5712_ (.A(net58),
    .Y(_4080_));
 sky130_fd_sc_hs__inv_1 _5713_ (.A(net59),
    .Y(_4086_));
 sky130_fd_sc_hs__inv_1 _5714_ (.A(net60),
    .Y(_4092_));
 sky130_fd_sc_hs__inv_1 _5715_ (.A(net61),
    .Y(_4098_));
 sky130_fd_sc_hs__inv_1 _5716_ (.A(net62),
    .Y(_4104_));
 sky130_fd_sc_hs__inv_1 _5717_ (.A(net63),
    .Y(_4110_));
 sky130_fd_sc_hs__inv_1 _5718_ (.A(net65),
    .Y(_4116_));
 sky130_fd_sc_hs__inv_1 _5719_ (.A(_3732_),
    .Y(_2288_));
 sky130_fd_sc_hs__inv_1 _5720_ (.A(_3744_),
    .Y(_2306_));
 sky130_fd_sc_hs__inv_1 _5721_ (.A(_3758_),
    .Y(_2373_));
 sky130_fd_sc_hs__inv_1 _5722_ (.A(_3772_),
    .Y(_2401_));
 sky130_fd_sc_hs__inv_1 _5723_ (.A(_3780_),
    .Y(_2440_));
 sky130_fd_sc_hs__inv_1 _5724_ (.A(_3810_),
    .Y(_2642_));
 sky130_fd_sc_hs__inv_1 _5725_ (.A(_3820_),
    .Y(_2696_));
 sky130_fd_sc_hs__inv_1 _5726_ (.A(_3721_),
    .Y(_2250_));
 sky130_fd_sc_hs__inv_1 _5727_ (.A(_3796_),
    .Y(_2523_));
 sky130_fd_sc_hs__inv_1 _5728_ (.A(_3830_),
    .Y(_2831_));
 sky130_fd_sc_hs__mux2_1 _5729_ (.A0(\genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0] ),
    .A1(\genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[2] ),
    .S(_0088_),
    .X(_0006_));
 sky130_fd_sc_hs__mux2_1 _5730_ (.A0(\genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[2] ),
    .A1(_0084_),
    .S(_0088_),
    .X(_0007_));
 sky130_fd_sc_hs__buf_8 _5731_ (.A(_0381_),
    .X(_0810_));
 sky130_fd_sc_hs__o21ai_4 _5732_ (.A1(_0092_),
    .A2(net187),
    .B1(net79),
    .Y(_0811_));
 sky130_fd_sc_hs__buf_8 _5733_ (.A(_0811_),
    .X(_0812_));
 sky130_fd_sc_hs__mux2i_1 _5734_ (.A0(_0392_),
    .A1(_0810_),
    .S(_0812_),
    .Y(_0008_));
 sky130_fd_sc_hs__inv_2 _5735_ (.A(_0090_),
    .Y(_0813_));
 sky130_fd_sc_hs__buf_8 _5736_ (.A(_0813_),
    .X(_0814_));
 sky130_fd_sc_hs__nand2_8 _5737_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .B(_0094_),
    .Y(_0815_));
 sky130_fd_sc_hs__buf_4 _5738_ (.A(_0815_),
    .X(_0816_));
 sky130_fd_sc_hs__o21ai_1 _5739_ (.A1(_0814_),
    .A2(_0094_),
    .B1(_0816_),
    .Y(_0009_));
 sky130_fd_sc_hs__nand2_1 _5740_ (.A(_0123_),
    .B(_0812_),
    .Y(_0817_));
 sky130_fd_sc_hs__o21ai_1 _5741_ (.A1(_0092_),
    .A2(_0812_),
    .B1(_0817_),
    .Y(_0010_));
 sky130_fd_sc_hs__nor2b_4 _5742_ (.A(net185),
    .B_N(net186),
    .Y(_0818_));
 sky130_fd_sc_hs__nand2_8 _5743_ (.A(_0122_),
    .B(_0818_),
    .Y(_0819_));
 sky130_fd_sc_hs__nor2_1 _5744_ (.A(_0812_),
    .B(_0819_),
    .Y(_0820_));
 sky130_fd_sc_hs__mux2_1 _5745_ (.A0(\genblk3.gen_multdiv_fast.multdiv_i.div_by_zero_q ),
    .A1(_0531_),
    .S(_0820_),
    .X(_0011_));
 sky130_fd_sc_hs__nor4_4 _5746_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.md_state_q[2] ),
    .B(\genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .C(_0122_),
    .D(_0811_),
    .Y(_0821_));
 sky130_fd_sc_hs__nor2_1 _5747_ (.A(_0590_),
    .B(_0094_),
    .Y(_0822_));
 sky130_fd_sc_hs__a21oi_1 _5748_ (.A1(_0590_),
    .A2(_0821_),
    .B1(_0822_),
    .Y(_0012_));
 sky130_fd_sc_hs__clkbuf_8 _5749_ (.A(_3705_),
    .X(_0823_));
 sky130_fd_sc_hs__a22oi_1 _5750_ (.A1(_3703_),
    .A2(_0812_),
    .B1(_0821_),
    .B2(_0823_),
    .Y(_0013_));
 sky130_fd_sc_hs__nand2b_1 _5751_ (.A_N(_3706_),
    .B(_0821_),
    .Y(_0824_));
 sky130_fd_sc_hs__a21oi_1 _5752_ (.A1(_0094_),
    .A2(_0824_),
    .B1(_0098_),
    .Y(_0825_));
 sky130_fd_sc_hs__a31oi_1 _5753_ (.A1(_0098_),
    .A2(_3706_),
    .A3(_0821_),
    .B1(_0825_),
    .Y(_0014_));
 sky130_fd_sc_hs__clkinv_4 _5754_ (.A(_0097_),
    .Y(_0826_));
 sky130_fd_sc_hs__nor3_4 _5755_ (.A(_0098_),
    .B(_0590_),
    .C(\genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .Y(_0827_));
 sky130_fd_sc_hs__xnor2_4 _5756_ (.A(_0097_),
    .B(_0827_),
    .Y(_0828_));
 sky130_fd_sc_hs__a22oi_1 _5757_ (.A1(_0826_),
    .A2(_0812_),
    .B1(_0821_),
    .B2(_0828_),
    .Y(_0015_));
 sky130_fd_sc_hs__nor3b_4 _5758_ (.A(_0097_),
    .B(_0098_),
    .C_N(_3706_),
    .Y(_0829_));
 sky130_fd_sc_hs__nand2b_1 _5759_ (.A_N(_0829_),
    .B(_0821_),
    .Y(_0830_));
 sky130_fd_sc_hs__a21oi_1 _5760_ (.A1(_0094_),
    .A2(_0830_),
    .B1(_0096_),
    .Y(_0831_));
 sky130_fd_sc_hs__a31oi_1 _5761_ (.A1(_0096_),
    .A2(_0821_),
    .A3(_0829_),
    .B1(_0831_),
    .Y(_0016_));
 sky130_fd_sc_hs__nor2_2 _5762_ (.A(_0383_),
    .B(_0812_),
    .Y(_0832_));
 sky130_fd_sc_hs__clkbuf_8 _5763_ (.A(_0832_),
    .X(_0833_));
 sky130_fd_sc_hs__clkbuf_4 _5764_ (.A(_0833_),
    .X(_0834_));
 sky130_fd_sc_hs__clkbuf_16 _5765_ (.A(_0513_),
    .X(_0835_));
 sky130_fd_sc_hs__buf_8 _5766_ (.A(_0835_),
    .X(_0836_));
 sky130_fd_sc_hs__mux2i_4 _5767_ (.A0(net121),
    .A1(net191),
    .S(_0836_),
    .Y(_0837_));
 sky130_fd_sc_hs__clkbuf_4 _5768_ (.A(_0832_),
    .X(_0838_));
 sky130_fd_sc_hs__nor2_1 _5769_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[0] ),
    .B(_0838_),
    .Y(_0839_));
 sky130_fd_sc_hs__a21oi_1 _5770_ (.A1(_0834_),
    .A2(_0837_),
    .B1(_0839_),
    .Y(_0017_));
 sky130_fd_sc_hs__nor2_1 _5771_ (.A(net122),
    .B(_0836_),
    .Y(_0840_));
 sky130_fd_sc_hs__nand2_8 _5772_ (.A(net145),
    .B(net188),
    .Y(_0841_));
 sky130_fd_sc_hs__clkbuf_8 _5773_ (.A(_0841_),
    .X(_0842_));
 sky130_fd_sc_hs__nor2_1 _5774_ (.A(net192),
    .B(_0842_),
    .Y(_0843_));
 sky130_fd_sc_hs__nand2_1 _5775_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[10] ),
    .B(_0816_),
    .Y(_0844_));
 sky130_fd_sc_hs__o31ai_1 _5776_ (.A1(_0815_),
    .A2(_0840_),
    .A3(_0843_),
    .B1(_0844_),
    .Y(_0018_));
 sky130_fd_sc_hs__mux2i_4 _5777_ (.A0(net123),
    .A1(net193),
    .S(_0836_),
    .Y(_0845_));
 sky130_fd_sc_hs__nor2_1 _5778_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[11] ),
    .B(_0838_),
    .Y(_0846_));
 sky130_fd_sc_hs__a21oi_1 _5779_ (.A1(_0834_),
    .A2(_0845_),
    .B1(_0846_),
    .Y(_0019_));
 sky130_fd_sc_hs__nor3_4 _5780_ (.A(_0333_),
    .B(_0335_),
    .C(_0841_),
    .Y(_0847_));
 sky130_fd_sc_hs__a21oi_4 _5781_ (.A1(net124),
    .A2(_0842_),
    .B1(_0847_),
    .Y(_0848_));
 sky130_fd_sc_hs__nor2_1 _5782_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[12] ),
    .B(_0838_),
    .Y(_0849_));
 sky130_fd_sc_hs__a21oi_1 _5783_ (.A1(_0834_),
    .A2(_0848_),
    .B1(_0849_),
    .Y(_0020_));
 sky130_fd_sc_hs__mux2i_4 _5784_ (.A0(net125),
    .A1(net195),
    .S(_0836_),
    .Y(_0850_));
 sky130_fd_sc_hs__nor2_1 _5785_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[13] ),
    .B(_0838_),
    .Y(_0851_));
 sky130_fd_sc_hs__a21oi_1 _5786_ (.A1(_0834_),
    .A2(_0850_),
    .B1(_0851_),
    .Y(_0021_));
 sky130_fd_sc_hs__mux2i_4 _5787_ (.A0(net126),
    .A1(net16),
    .S(_0836_),
    .Y(_0852_));
 sky130_fd_sc_hs__nor2_1 _5788_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[14] ),
    .B(_0838_),
    .Y(_0853_));
 sky130_fd_sc_hs__a21oi_1 _5789_ (.A1(_0834_),
    .A2(_0852_),
    .B1(_0853_),
    .Y(_0022_));
 sky130_fd_sc_hs__buf_16 _5790_ (.A(_0835_),
    .X(_0854_));
 sky130_fd_sc_hs__mux2i_4 _5791_ (.A0(net127),
    .A1(net15),
    .S(_0854_),
    .Y(_0855_));
 sky130_fd_sc_hs__nor2_1 _5792_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[15] ),
    .B(_0838_),
    .Y(_0856_));
 sky130_fd_sc_hs__a21oi_1 _5793_ (.A1(_0834_),
    .A2(_0855_),
    .B1(_0856_),
    .Y(_0023_));
 sky130_fd_sc_hs__mux2i_4 _5794_ (.A0(net128),
    .A1(net198),
    .S(_0854_),
    .Y(_0857_));
 sky130_fd_sc_hs__nor2_1 _5795_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[16] ),
    .B(_0838_),
    .Y(_0858_));
 sky130_fd_sc_hs__a21oi_1 _5796_ (.A1(_0834_),
    .A2(_0857_),
    .B1(_0858_),
    .Y(_0024_));
 sky130_fd_sc_hs__mux2i_4 _5797_ (.A0(net129),
    .A1(net199),
    .S(_0854_),
    .Y(_0859_));
 sky130_fd_sc_hs__clkbuf_4 _5798_ (.A(_0832_),
    .X(_0860_));
 sky130_fd_sc_hs__nor2_1 _5799_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[17] ),
    .B(_0860_),
    .Y(_0861_));
 sky130_fd_sc_hs__a21oi_1 _5800_ (.A1(_0834_),
    .A2(_0859_),
    .B1(_0861_),
    .Y(_0025_));
 sky130_fd_sc_hs__mux2i_4 _5801_ (.A0(net130),
    .A1(net200),
    .S(_0854_),
    .Y(_0862_));
 sky130_fd_sc_hs__nor2_1 _5802_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[18] ),
    .B(_0860_),
    .Y(_0863_));
 sky130_fd_sc_hs__a21oi_1 _5803_ (.A1(_0834_),
    .A2(_0862_),
    .B1(_0863_),
    .Y(_0026_));
 sky130_fd_sc_hs__mux2i_4 _5804_ (.A0(net131),
    .A1(net201),
    .S(_0854_),
    .Y(_0864_));
 sky130_fd_sc_hs__nor2_1 _5805_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[19] ),
    .B(_0860_),
    .Y(_0865_));
 sky130_fd_sc_hs__a21oi_1 _5806_ (.A1(_0834_),
    .A2(_0864_),
    .B1(_0865_),
    .Y(_0027_));
 sky130_fd_sc_hs__nor2_1 _5807_ (.A(_0306_),
    .B(_0841_),
    .Y(_0866_));
 sky130_fd_sc_hs__a21oi_4 _5808_ (.A1(net132),
    .A2(_0842_),
    .B1(_0866_),
    .Y(_0867_));
 sky130_fd_sc_hs__nand2_1 _5809_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[1] ),
    .B(_0816_),
    .Y(_0868_));
 sky130_fd_sc_hs__o21ai_1 _5810_ (.A1(_0816_),
    .A2(_0867_),
    .B1(_0868_),
    .Y(_0028_));
 sky130_fd_sc_hs__nor2_1 _5811_ (.A(net133),
    .B(_0836_),
    .Y(_0869_));
 sky130_fd_sc_hs__nor2_1 _5812_ (.A(net203),
    .B(_0842_),
    .Y(_0870_));
 sky130_fd_sc_hs__nand2_1 _5813_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[20] ),
    .B(_0816_),
    .Y(_0871_));
 sky130_fd_sc_hs__o31ai_1 _5814_ (.A1(_0815_),
    .A2(_0869_),
    .A3(_0870_),
    .B1(_0871_),
    .Y(_0029_));
 sky130_fd_sc_hs__clkbuf_4 _5815_ (.A(_0833_),
    .X(_0872_));
 sky130_fd_sc_hs__mux2i_2 _5816_ (.A0(net134),
    .A1(net204),
    .S(_0854_),
    .Y(_0873_));
 sky130_fd_sc_hs__nor2_1 _5817_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[21] ),
    .B(_0860_),
    .Y(_0874_));
 sky130_fd_sc_hs__a21oi_1 _5818_ (.A1(_0872_),
    .A2(_0873_),
    .B1(_0874_),
    .Y(_0030_));
 sky130_fd_sc_hs__mux2i_4 _5819_ (.A0(net135),
    .A1(net205),
    .S(_0854_),
    .Y(_0875_));
 sky130_fd_sc_hs__nor2_1 _5820_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[22] ),
    .B(_0860_),
    .Y(_0876_));
 sky130_fd_sc_hs__a21oi_1 _5821_ (.A1(_0872_),
    .A2(_0875_),
    .B1(_0876_),
    .Y(_0031_));
 sky130_fd_sc_hs__mux2i_2 _5822_ (.A0(net136),
    .A1(net206),
    .S(_0854_),
    .Y(_0877_));
 sky130_fd_sc_hs__nor2_1 _5823_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[23] ),
    .B(_0860_),
    .Y(_0878_));
 sky130_fd_sc_hs__a21oi_1 _5824_ (.A1(_0872_),
    .A2(_0877_),
    .B1(_0878_),
    .Y(_0032_));
 sky130_fd_sc_hs__mux2i_4 _5825_ (.A0(net137),
    .A1(net13),
    .S(_0854_),
    .Y(_0879_));
 sky130_fd_sc_hs__nor2_1 _5826_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[24] ),
    .B(_0860_),
    .Y(_0880_));
 sky130_fd_sc_hs__a21oi_1 _5827_ (.A1(_0872_),
    .A2(_0879_),
    .B1(_0880_),
    .Y(_0033_));
 sky130_fd_sc_hs__mux2i_4 _5828_ (.A0(net138),
    .A1(net208),
    .S(_0854_),
    .Y(_0881_));
 sky130_fd_sc_hs__nor2_1 _5829_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[25] ),
    .B(_0860_),
    .Y(_0882_));
 sky130_fd_sc_hs__a21oi_1 _5830_ (.A1(_0872_),
    .A2(_0881_),
    .B1(_0882_),
    .Y(_0034_));
 sky130_fd_sc_hs__mux2i_4 _5831_ (.A0(net139),
    .A1(net209),
    .S(_0835_),
    .Y(_0883_));
 sky130_fd_sc_hs__nor2_1 _5832_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[26] ),
    .B(_0860_),
    .Y(_0884_));
 sky130_fd_sc_hs__a21oi_1 _5833_ (.A1(_0872_),
    .A2(_0883_),
    .B1(_0884_),
    .Y(_0035_));
 sky130_fd_sc_hs__nor2_1 _5834_ (.A(net140),
    .B(_0836_),
    .Y(_0885_));
 sky130_fd_sc_hs__nor2_1 _5835_ (.A(net210),
    .B(_0842_),
    .Y(_0886_));
 sky130_fd_sc_hs__nand2_1 _5836_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[27] ),
    .B(_0816_),
    .Y(_0887_));
 sky130_fd_sc_hs__o31ai_1 _5837_ (.A1(_0815_),
    .A2(_0885_),
    .A3(_0886_),
    .B1(_0887_),
    .Y(_0036_));
 sky130_fd_sc_hs__mux2i_2 _5838_ (.A0(net141),
    .A1(net12),
    .S(_0835_),
    .Y(_0888_));
 sky130_fd_sc_hs__nor2_1 _5839_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[28] ),
    .B(_0860_),
    .Y(_0889_));
 sky130_fd_sc_hs__a21oi_1 _5840_ (.A1(_0872_),
    .A2(_0888_),
    .B1(_0889_),
    .Y(_0037_));
 sky130_fd_sc_hs__mux2i_2 _5841_ (.A0(net142),
    .A1(net9),
    .S(_0835_),
    .Y(_0890_));
 sky130_fd_sc_hs__nor2_1 _5842_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[29] ),
    .B(_0833_),
    .Y(_0891_));
 sky130_fd_sc_hs__a21oi_1 _5843_ (.A1(_0872_),
    .A2(_0890_),
    .B1(_0891_),
    .Y(_0038_));
 sky130_fd_sc_hs__mux2i_4 _5844_ (.A0(net143),
    .A1(net213),
    .S(_0835_),
    .Y(_0892_));
 sky130_fd_sc_hs__nor2_1 _5845_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[2] ),
    .B(_0833_),
    .Y(_0893_));
 sky130_fd_sc_hs__a21oi_1 _5846_ (.A1(_0872_),
    .A2(_0892_),
    .B1(_0893_),
    .Y(_0039_));
 sky130_fd_sc_hs__nor2_1 _5847_ (.A(net144),
    .B(_0836_),
    .Y(_0894_));
 sky130_fd_sc_hs__nor2_1 _5848_ (.A(net214),
    .B(_0842_),
    .Y(_0895_));
 sky130_fd_sc_hs__nand2_1 _5849_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[30] ),
    .B(_0816_),
    .Y(_0896_));
 sky130_fd_sc_hs__o31ai_1 _5850_ (.A1(_0815_),
    .A2(_0894_),
    .A3(_0895_),
    .B1(_0896_),
    .Y(_0040_));
 sky130_fd_sc_hs__nand2_1 _5851_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[31] ),
    .B(_0816_),
    .Y(_0897_));
 sky130_fd_sc_hs__o211ai_1 _5852_ (.A1(_0522_),
    .A2(net215),
    .B1(_0833_),
    .C1(net145),
    .Y(_0898_));
 sky130_fd_sc_hs__nand2_1 _5853_ (.A(_0897_),
    .B(_0898_),
    .Y(_0041_));
 sky130_fd_sc_hs__mux2i_4 _5854_ (.A0(net146),
    .A1(net216),
    .S(_0835_),
    .Y(_0899_));
 sky130_fd_sc_hs__nor2_1 _5855_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[3] ),
    .B(_0833_),
    .Y(_0900_));
 sky130_fd_sc_hs__a21oi_1 _5856_ (.A1(_0872_),
    .A2(_0899_),
    .B1(_0900_),
    .Y(_0042_));
 sky130_fd_sc_hs__nor2_1 _5857_ (.A(net147),
    .B(_0836_),
    .Y(_0901_));
 sky130_fd_sc_hs__nor2_1 _5858_ (.A(net217),
    .B(_0842_),
    .Y(_0902_));
 sky130_fd_sc_hs__nand2_1 _5859_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[4] ),
    .B(_0815_),
    .Y(_0903_));
 sky130_fd_sc_hs__o31ai_1 _5860_ (.A1(_0815_),
    .A2(_0901_),
    .A3(_0902_),
    .B1(_0903_),
    .Y(_0043_));
 sky130_fd_sc_hs__nor2_1 _5861_ (.A(_0317_),
    .B(_0841_),
    .Y(_0904_));
 sky130_fd_sc_hs__a21oi_4 _5862_ (.A1(net148),
    .A2(_0842_),
    .B1(_0904_),
    .Y(_0905_));
 sky130_fd_sc_hs__nor2_1 _5863_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[5] ),
    .B(_0833_),
    .Y(_0906_));
 sky130_fd_sc_hs__a21oi_1 _5864_ (.A1(_0838_),
    .A2(_0905_),
    .B1(_0906_),
    .Y(_0044_));
 sky130_fd_sc_hs__mux2i_4 _5865_ (.A0(net149),
    .A1(net219),
    .S(_0835_),
    .Y(_0907_));
 sky130_fd_sc_hs__nor2_1 _5866_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[6] ),
    .B(_0833_),
    .Y(_0908_));
 sky130_fd_sc_hs__a21oi_1 _5867_ (.A1(_0838_),
    .A2(_0907_),
    .B1(_0908_),
    .Y(_0045_));
 sky130_fd_sc_hs__mux2i_4 _5868_ (.A0(net150),
    .A1(net220),
    .S(_0835_),
    .Y(_0909_));
 sky130_fd_sc_hs__nor2_1 _5869_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[7] ),
    .B(_0833_),
    .Y(_0910_));
 sky130_fd_sc_hs__a21oi_1 _5870_ (.A1(_0838_),
    .A2(_0909_),
    .B1(_0910_),
    .Y(_0046_));
 sky130_fd_sc_hs__nor2_1 _5871_ (.A(net151),
    .B(_0836_),
    .Y(_0911_));
 sky130_fd_sc_hs__nor2_1 _5872_ (.A(net221),
    .B(_0842_),
    .Y(_0912_));
 sky130_fd_sc_hs__nand2_1 _5873_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[8] ),
    .B(_0815_),
    .Y(_0913_));
 sky130_fd_sc_hs__o31ai_1 _5874_ (.A1(_0815_),
    .A2(_0911_),
    .A3(_0912_),
    .B1(_0913_),
    .Y(_0047_));
 sky130_fd_sc_hs__nor2_1 _5875_ (.A(_0299_),
    .B(_0841_),
    .Y(_0914_));
 sky130_fd_sc_hs__a21oi_1 _5876_ (.A1(net152),
    .A2(_0842_),
    .B1(_0914_),
    .Y(_0915_));
 sky130_fd_sc_hs__nand2_1 _5877_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[9] ),
    .B(_0816_),
    .Y(_0916_));
 sky130_fd_sc_hs__o21ai_1 _5878_ (.A1(_0816_),
    .A2(_0915_),
    .B1(_0916_),
    .Y(_0048_));
 sky130_fd_sc_hs__nor2_8 _5879_ (.A(_0102_),
    .B(_0815_),
    .Y(_0917_));
 sky130_fd_sc_hs__buf_4 _5880_ (.A(_0917_),
    .X(_0918_));
 sky130_fd_sc_hs__nor2_1 _5881_ (.A(_0096_),
    .B(_0098_),
    .Y(_0919_));
 sky130_fd_sc_hs__buf_8 _5882_ (.A(_3704_),
    .X(_0920_));
 sky130_fd_sc_hs__nor2_4 _5883_ (.A(_0391_),
    .B(_0812_),
    .Y(_0921_));
 sky130_fd_sc_hs__and2_2 _5884_ (.A(_0920_),
    .B(_0921_),
    .X(_0922_));
 sky130_fd_sc_hs__o21a_1 _5885_ (.A1(_0265_),
    .A2(_0270_),
    .B1(_0275_),
    .X(_0923_));
 sky130_fd_sc_hs__nand2_1 _5886_ (.A(_0401_),
    .B(_0402_),
    .Y(_0924_));
 sky130_fd_sc_hs__nor2_1 _5887_ (.A(net105),
    .B(_0407_),
    .Y(_0925_));
 sky130_fd_sc_hs__nor2_1 _5888_ (.A(_0385_),
    .B(_0407_),
    .Y(_0926_));
 sky130_fd_sc_hs__o221ai_2 _5889_ (.A1(_0923_),
    .A2(_0924_),
    .B1(_0925_),
    .B2(_0926_),
    .C1(_0400_),
    .Y(_0927_));
 sky130_fd_sc_hs__a2111o_1 _5890_ (.A1(_0385_),
    .A2(net105),
    .B1(_0923_),
    .C1(_0400_),
    .D1(_0924_),
    .X(_0928_));
 sky130_fd_sc_hs__o221ai_1 _5891_ (.A1(_0382_),
    .A2(_0390_),
    .B1(_0395_),
    .B2(_0399_),
    .C1(_0407_),
    .Y(_0929_));
 sky130_fd_sc_hs__o21a_1 _5892_ (.A1(_0385_),
    .A2(net105),
    .B1(_0929_),
    .X(_0930_));
 sky130_fd_sc_hs__and3_4 _5893_ (.A(_0927_),
    .B(_0928_),
    .C(_0930_),
    .X(_0931_));
 sky130_fd_sc_hs__buf_8 _5894_ (.A(_0931_),
    .X(_0932_));
 sky130_fd_sc_hs__nor2_8 _5895_ (.A(_0097_),
    .B(_0932_),
    .Y(_0933_));
 sky130_fd_sc_hs__and2_1 _5896_ (.A(_0922_),
    .B(_0933_),
    .X(_0934_));
 sky130_fd_sc_hs__a21oi_1 _5897_ (.A1(_0919_),
    .A2(_0934_),
    .B1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[0] ),
    .Y(_0935_));
 sky130_fd_sc_hs__nor2_1 _5898_ (.A(_0918_),
    .B(_0935_),
    .Y(_0049_));
 sky130_fd_sc_hs__clkinv_2 _5899_ (.A(_0919_),
    .Y(_0936_));
 sky130_fd_sc_hs__nor3_4 _5900_ (.A(_0826_),
    .B(_0936_),
    .C(_0932_),
    .Y(_0937_));
 sky130_fd_sc_hs__buf_8 _5901_ (.A(_3708_),
    .X(_0938_));
 sky130_fd_sc_hs__and2_4 _5902_ (.A(_0938_),
    .B(_0921_),
    .X(_0939_));
 sky130_fd_sc_hs__a21oi_1 _5903_ (.A1(_0937_),
    .A2(_0939_),
    .B1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[10] ),
    .Y(_0940_));
 sky130_fd_sc_hs__nor2_1 _5904_ (.A(_0918_),
    .B(_0940_),
    .Y(_0050_));
 sky130_fd_sc_hs__buf_8 _5905_ (.A(_3712_),
    .X(_0941_));
 sky130_fd_sc_hs__and2_4 _5906_ (.A(_0941_),
    .B(_0921_),
    .X(_0942_));
 sky130_fd_sc_hs__a21oi_1 _5907_ (.A1(_0937_),
    .A2(_0942_),
    .B1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[11] ),
    .Y(_0943_));
 sky130_fd_sc_hs__nor2_1 _5908_ (.A(_0918_),
    .B(_0943_),
    .Y(_0051_));
 sky130_fd_sc_hs__nand2b_2 _5909_ (.A_N(_0096_),
    .B(_0098_),
    .Y(_0944_));
 sky130_fd_sc_hs__nor3_4 _5910_ (.A(_0826_),
    .B(_0931_),
    .C(_0944_),
    .Y(_0945_));
 sky130_fd_sc_hs__a21oi_1 _5911_ (.A1(_0922_),
    .A2(_0945_),
    .B1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[12] ),
    .Y(_0946_));
 sky130_fd_sc_hs__nor2_1 _5912_ (.A(_0918_),
    .B(_0946_),
    .Y(_0052_));
 sky130_fd_sc_hs__and2_4 _5913_ (.A(_0095_),
    .B(_0921_),
    .X(_0947_));
 sky130_fd_sc_hs__a21oi_1 _5914_ (.A1(_0945_),
    .A2(_0947_),
    .B1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[13] ),
    .Y(_0948_));
 sky130_fd_sc_hs__nor2_1 _5915_ (.A(_0918_),
    .B(_0948_),
    .Y(_0053_));
 sky130_fd_sc_hs__a21oi_1 _5916_ (.A1(_0939_),
    .A2(_0945_),
    .B1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[14] ),
    .Y(_0949_));
 sky130_fd_sc_hs__nor2_1 _5917_ (.A(_0918_),
    .B(_0949_),
    .Y(_0054_));
 sky130_fd_sc_hs__a21oi_1 _5918_ (.A1(_0942_),
    .A2(_0945_),
    .B1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[15] ),
    .Y(_0950_));
 sky130_fd_sc_hs__nor2_1 _5919_ (.A(_0918_),
    .B(_0950_),
    .Y(_0055_));
 sky130_fd_sc_hs__nor2b_4 _5920_ (.A(_0098_),
    .B_N(_0096_),
    .Y(_0951_));
 sky130_fd_sc_hs__a21oi_1 _5921_ (.A1(_0934_),
    .A2(_0951_),
    .B1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[16] ),
    .Y(_0952_));
 sky130_fd_sc_hs__nor2_1 _5922_ (.A(_0918_),
    .B(_0952_),
    .Y(_0056_));
 sky130_fd_sc_hs__nand2_4 _5923_ (.A(_0433_),
    .B(_0833_),
    .Y(_0953_));
 sky130_fd_sc_hs__and2_2 _5924_ (.A(_0933_),
    .B(_0951_),
    .X(_0954_));
 sky130_fd_sc_hs__a22o_1 _5925_ (.A1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[17] ),
    .A2(_0953_),
    .B1(_0947_),
    .B2(_0954_),
    .X(_0057_));
 sky130_fd_sc_hs__a21oi_1 _5926_ (.A1(_0939_),
    .A2(_0954_),
    .B1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[18] ),
    .Y(_0955_));
 sky130_fd_sc_hs__nor2_1 _5927_ (.A(_0918_),
    .B(_0955_),
    .Y(_0058_));
 sky130_fd_sc_hs__a21oi_1 _5928_ (.A1(_0942_),
    .A2(_0954_),
    .B1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[19] ),
    .Y(_0956_));
 sky130_fd_sc_hs__nor2_1 _5929_ (.A(_0918_),
    .B(_0956_),
    .Y(_0059_));
 sky130_fd_sc_hs__nand3_1 _5930_ (.A(_0927_),
    .B(_0928_),
    .C(_0930_),
    .Y(_0957_));
 sky130_fd_sc_hs__buf_8 _5931_ (.A(_0957_),
    .X(_0958_));
 sky130_fd_sc_hs__buf_8 _5932_ (.A(_0958_),
    .X(_0959_));
 sky130_fd_sc_hs__a32o_1 _5933_ (.A1(_0100_),
    .A2(_0921_),
    .A3(_0959_),
    .B1(_0953_),
    .B2(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[1] ),
    .X(_0060_));
 sky130_fd_sc_hs__buf_4 _5934_ (.A(_0917_),
    .X(_0960_));
 sky130_fd_sc_hs__and2_1 _5935_ (.A(_0096_),
    .B(_0098_),
    .X(_0961_));
 sky130_fd_sc_hs__buf_4 _5936_ (.A(_0961_),
    .X(_0962_));
 sky130_fd_sc_hs__a21oi_1 _5937_ (.A1(_0934_),
    .A2(_0962_),
    .B1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[20] ),
    .Y(_0963_));
 sky130_fd_sc_hs__nor2_1 _5938_ (.A(_0960_),
    .B(_0963_),
    .Y(_0061_));
 sky130_fd_sc_hs__and2_2 _5939_ (.A(_0933_),
    .B(_0962_),
    .X(_0964_));
 sky130_fd_sc_hs__a21oi_1 _5940_ (.A1(_0947_),
    .A2(_0964_),
    .B1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[21] ),
    .Y(_0965_));
 sky130_fd_sc_hs__nor2_1 _5941_ (.A(_0960_),
    .B(_0965_),
    .Y(_0062_));
 sky130_fd_sc_hs__a21oi_1 _5942_ (.A1(_0939_),
    .A2(_0964_),
    .B1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[22] ),
    .Y(_0966_));
 sky130_fd_sc_hs__nor2_1 _5943_ (.A(_0960_),
    .B(_0966_),
    .Y(_0063_));
 sky130_fd_sc_hs__a21oi_1 _5944_ (.A1(_0942_),
    .A2(_0964_),
    .B1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[23] ),
    .Y(_0967_));
 sky130_fd_sc_hs__nor2_1 _5945_ (.A(_0960_),
    .B(_0967_),
    .Y(_0064_));
 sky130_fd_sc_hs__and3_1 _5946_ (.A(_0097_),
    .B(_0958_),
    .C(_0951_),
    .X(_0968_));
 sky130_fd_sc_hs__clkbuf_4 _5947_ (.A(_0968_),
    .X(_0969_));
 sky130_fd_sc_hs__a21oi_1 _5948_ (.A1(_0922_),
    .A2(_0969_),
    .B1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[24] ),
    .Y(_0970_));
 sky130_fd_sc_hs__nor2_1 _5949_ (.A(_0960_),
    .B(_0970_),
    .Y(_0065_));
 sky130_fd_sc_hs__a21oi_1 _5950_ (.A1(_0947_),
    .A2(_0969_),
    .B1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[25] ),
    .Y(_0971_));
 sky130_fd_sc_hs__nor2_1 _5951_ (.A(_0960_),
    .B(_0971_),
    .Y(_0066_));
 sky130_fd_sc_hs__a21oi_1 _5952_ (.A1(_0939_),
    .A2(_0969_),
    .B1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[26] ),
    .Y(_0972_));
 sky130_fd_sc_hs__nor2_1 _5953_ (.A(_0960_),
    .B(_0972_),
    .Y(_0067_));
 sky130_fd_sc_hs__a21oi_1 _5954_ (.A1(_0942_),
    .A2(_0969_),
    .B1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[27] ),
    .Y(_0973_));
 sky130_fd_sc_hs__nor2_1 _5955_ (.A(_0960_),
    .B(_0973_),
    .Y(_0068_));
 sky130_fd_sc_hs__nor2_2 _5956_ (.A(_0826_),
    .B(_0932_),
    .Y(_0974_));
 sky130_fd_sc_hs__and2_2 _5957_ (.A(_0974_),
    .B(_0962_),
    .X(_0975_));
 sky130_fd_sc_hs__a22o_1 _5958_ (.A1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[28] ),
    .A2(_0953_),
    .B1(_0922_),
    .B2(_0975_),
    .X(_0069_));
 sky130_fd_sc_hs__a21oi_1 _5959_ (.A1(_0947_),
    .A2(_0975_),
    .B1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[29] ),
    .Y(_0976_));
 sky130_fd_sc_hs__nor2_1 _5960_ (.A(_0960_),
    .B(_0976_),
    .Y(_0070_));
 sky130_fd_sc_hs__nor3_4 _5961_ (.A(_0097_),
    .B(_0936_),
    .C(_0932_),
    .Y(_0977_));
 sky130_fd_sc_hs__a21oi_1 _5962_ (.A1(_0939_),
    .A2(_0977_),
    .B1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[2] ),
    .Y(_0978_));
 sky130_fd_sc_hs__nor2_1 _5963_ (.A(_0960_),
    .B(_0978_),
    .Y(_0071_));
 sky130_fd_sc_hs__a21oi_1 _5964_ (.A1(_0939_),
    .A2(_0975_),
    .B1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[30] ),
    .Y(_0979_));
 sky130_fd_sc_hs__nor2_1 _5965_ (.A(_0917_),
    .B(_0979_),
    .Y(_0072_));
 sky130_fd_sc_hs__a21oi_1 _5966_ (.A1(_0942_),
    .A2(_0975_),
    .B1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[31] ),
    .Y(_0980_));
 sky130_fd_sc_hs__nor2_1 _5967_ (.A(_0917_),
    .B(_0980_),
    .Y(_0073_));
 sky130_fd_sc_hs__a21oi_1 _5968_ (.A1(_0942_),
    .A2(_0977_),
    .B1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[3] ),
    .Y(_0981_));
 sky130_fd_sc_hs__nor2_1 _5969_ (.A(_0917_),
    .B(_0981_),
    .Y(_0074_));
 sky130_fd_sc_hs__nor2b_1 _5970_ (.A(_0096_),
    .B_N(_0098_),
    .Y(_0982_));
 sky130_fd_sc_hs__a21oi_1 _5971_ (.A1(_0934_),
    .A2(_0982_),
    .B1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[4] ),
    .Y(_0983_));
 sky130_fd_sc_hs__nor2_1 _5972_ (.A(_0917_),
    .B(_0983_),
    .Y(_0075_));
 sky130_fd_sc_hs__nor3_4 _5973_ (.A(_0097_),
    .B(_0932_),
    .C(_0944_),
    .Y(_0984_));
 sky130_fd_sc_hs__a21oi_1 _5974_ (.A1(_0947_),
    .A2(_0984_),
    .B1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[5] ),
    .Y(_0985_));
 sky130_fd_sc_hs__nor2_1 _5975_ (.A(_0917_),
    .B(_0985_),
    .Y(_0076_));
 sky130_fd_sc_hs__a21oi_1 _5976_ (.A1(_0939_),
    .A2(_0984_),
    .B1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[6] ),
    .Y(_0986_));
 sky130_fd_sc_hs__nor2_1 _5977_ (.A(_0917_),
    .B(_0986_),
    .Y(_0077_));
 sky130_fd_sc_hs__a21oi_1 _5978_ (.A1(_0942_),
    .A2(_0984_),
    .B1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[7] ),
    .Y(_0987_));
 sky130_fd_sc_hs__nor2_1 _5979_ (.A(_0917_),
    .B(_0987_),
    .Y(_0078_));
 sky130_fd_sc_hs__a21oi_1 _5980_ (.A1(_0922_),
    .A2(_0937_),
    .B1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[8] ),
    .Y(_0988_));
 sky130_fd_sc_hs__nor2_1 _5981_ (.A(_0917_),
    .B(_0988_),
    .Y(_0079_));
 sky130_fd_sc_hs__a22o_1 _5982_ (.A1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[9] ),
    .A2(_0953_),
    .B1(_0937_),
    .B2(_0947_),
    .X(_0080_));
 sky130_fd_sc_hs__nand3_4 _5983_ (.A(_0092_),
    .B(_0087_),
    .C(_0132_),
    .Y(net256));
 sky130_fd_sc_hs__buf_8 _5984_ (.A(_0517_),
    .X(_0989_));
 sky130_fd_sc_hs__buf_4 _5985_ (.A(_0989_),
    .X(_0990_));
 sky130_fd_sc_hs__nand2_1 _5986_ (.A(net191),
    .B(_0990_),
    .Y(_0991_));
 sky130_fd_sc_hs__nand2_8 _5987_ (.A(net177),
    .B(net189),
    .Y(_0992_));
 sky130_fd_sc_hs__buf_4 _5988_ (.A(_0992_),
    .X(_0993_));
 sky130_fd_sc_hs__nand2_1 _5989_ (.A(net153),
    .B(_0993_),
    .Y(_0994_));
 sky130_fd_sc_hs__clkbuf_4 _5990_ (.A(_0090_),
    .X(_0995_));
 sky130_fd_sc_hs__nor2_1 _5991_ (.A(_0995_),
    .B(net81),
    .Y(_0996_));
 sky130_fd_sc_hs__a311oi_4 _5992_ (.A1(_0091_),
    .A2(_0991_),
    .A3(_0994_),
    .B1(_0996_),
    .C1(_0788_),
    .Y(net257));
 sky130_fd_sc_hs__nor2_1 _5993_ (.A(net154),
    .B(_0989_),
    .Y(_0997_));
 sky130_fd_sc_hs__a311oi_1 _5994_ (.A1(_0341_),
    .A2(_0345_),
    .A3(_0989_),
    .B1(_0997_),
    .C1(_0813_),
    .Y(_0998_));
 sky130_fd_sc_hs__a21oi_2 _5995_ (.A1(_0814_),
    .A2(net82),
    .B1(_0998_),
    .Y(_0999_));
 sky130_fd_sc_hs__nor2_4 _5996_ (.A(_0109_),
    .B(_0999_),
    .Y(net258));
 sky130_fd_sc_hs__nand2_1 _5997_ (.A(net193),
    .B(_0990_),
    .Y(_1000_));
 sky130_fd_sc_hs__nand2_1 _5998_ (.A(net155),
    .B(_0993_),
    .Y(_1001_));
 sky130_fd_sc_hs__nor2_1 _5999_ (.A(_0995_),
    .B(net83),
    .Y(_1002_));
 sky130_fd_sc_hs__a311oi_4 _6000_ (.A1(_0091_),
    .A2(_1000_),
    .A3(_1001_),
    .B1(_1002_),
    .C1(_0788_),
    .Y(net259));
 sky130_fd_sc_hs__nand2_1 _6001_ (.A(net194),
    .B(_0990_),
    .Y(_1003_));
 sky130_fd_sc_hs__nand2_1 _6002_ (.A(net156),
    .B(_0993_),
    .Y(_1004_));
 sky130_fd_sc_hs__nor2_1 _6003_ (.A(_0995_),
    .B(net84),
    .Y(_1005_));
 sky130_fd_sc_hs__a311oi_4 _6004_ (.A1(_0091_),
    .A2(_1003_),
    .A3(_1004_),
    .B1(_1005_),
    .C1(_0788_),
    .Y(net260));
 sky130_fd_sc_hs__nand2_1 _6005_ (.A(net195),
    .B(_0990_),
    .Y(_1006_));
 sky130_fd_sc_hs__nand2_1 _6006_ (.A(net157),
    .B(_0993_),
    .Y(_1007_));
 sky130_fd_sc_hs__nor2_1 _6007_ (.A(_0995_),
    .B(net85),
    .Y(_1008_));
 sky130_fd_sc_hs__a311oi_4 _6008_ (.A1(_0091_),
    .A2(_1006_),
    .A3(_1007_),
    .B1(_1008_),
    .C1(_0788_),
    .Y(net261));
 sky130_fd_sc_hs__nand2_1 _6009_ (.A(net16),
    .B(_0990_),
    .Y(_1009_));
 sky130_fd_sc_hs__nand2_1 _6010_ (.A(net158),
    .B(_0993_),
    .Y(_1010_));
 sky130_fd_sc_hs__nor2_1 _6011_ (.A(_0995_),
    .B(net86),
    .Y(_1011_));
 sky130_fd_sc_hs__a311oi_4 _6012_ (.A1(_0091_),
    .A2(_1009_),
    .A3(_1010_),
    .B1(_1011_),
    .C1(_0788_),
    .Y(net262));
 sky130_fd_sc_hs__nand2_1 _6013_ (.A(net15),
    .B(_0990_),
    .Y(_1012_));
 sky130_fd_sc_hs__buf_4 _6014_ (.A(_0992_),
    .X(_1013_));
 sky130_fd_sc_hs__nand2_1 _6015_ (.A(net159),
    .B(_1013_),
    .Y(_1014_));
 sky130_fd_sc_hs__nor2_1 _6016_ (.A(_0995_),
    .B(net87),
    .Y(_1015_));
 sky130_fd_sc_hs__a311oi_4 _6017_ (.A1(_0091_),
    .A2(_1012_),
    .A3(_1014_),
    .B1(_1015_),
    .C1(_0788_),
    .Y(net263));
 sky130_fd_sc_hs__nand2_1 _6018_ (.A(net198),
    .B(_0990_),
    .Y(_1016_));
 sky130_fd_sc_hs__nand2_1 _6019_ (.A(net160),
    .B(_1013_),
    .Y(_1017_));
 sky130_fd_sc_hs__nor2_1 _6020_ (.A(_0995_),
    .B(net88),
    .Y(_1018_));
 sky130_fd_sc_hs__buf_8 _6021_ (.A(_0107_),
    .X(_1019_));
 sky130_fd_sc_hs__a311oi_4 _6022_ (.A1(_0091_),
    .A2(_1016_),
    .A3(_1017_),
    .B1(_1018_),
    .C1(_1019_),
    .Y(net264));
 sky130_fd_sc_hs__nand2_1 _6023_ (.A(net199),
    .B(_0990_),
    .Y(_1020_));
 sky130_fd_sc_hs__nand2_1 _6024_ (.A(net161),
    .B(_1013_),
    .Y(_1021_));
 sky130_fd_sc_hs__nor2_1 _6025_ (.A(_0995_),
    .B(net89),
    .Y(_1022_));
 sky130_fd_sc_hs__a311oi_4 _6026_ (.A1(_0091_),
    .A2(_1020_),
    .A3(_1021_),
    .B1(_1022_),
    .C1(_1019_),
    .Y(net265));
 sky130_fd_sc_hs__clkbuf_16 _6027_ (.A(_0090_),
    .X(_1023_));
 sky130_fd_sc_hs__nand2_1 _6028_ (.A(_0990_),
    .B(net200),
    .Y(_1024_));
 sky130_fd_sc_hs__nand2_1 _6029_ (.A(net162),
    .B(_1013_),
    .Y(_1025_));
 sky130_fd_sc_hs__nor2_1 _6030_ (.A(_0995_),
    .B(net90),
    .Y(_1026_));
 sky130_fd_sc_hs__a311oi_4 _6031_ (.A1(_1023_),
    .A2(_1024_),
    .A3(_1025_),
    .B1(_1026_),
    .C1(_1019_),
    .Y(net266));
 sky130_fd_sc_hs__nand2_1 _6032_ (.A(net201),
    .B(_0990_),
    .Y(_1027_));
 sky130_fd_sc_hs__nand2_1 _6033_ (.A(net163),
    .B(_1013_),
    .Y(_1028_));
 sky130_fd_sc_hs__buf_4 _6034_ (.A(_0090_),
    .X(_1029_));
 sky130_fd_sc_hs__nor2_1 _6035_ (.A(_1029_),
    .B(net91),
    .Y(_1030_));
 sky130_fd_sc_hs__a311oi_4 _6036_ (.A1(_1023_),
    .A2(_1027_),
    .A3(_1028_),
    .B1(_1030_),
    .C1(_1019_),
    .Y(net267));
 sky130_fd_sc_hs__nor2_1 _6037_ (.A(net164),
    .B(_0989_),
    .Y(_1031_));
 sky130_fd_sc_hs__a211oi_4 _6038_ (.A1(_0306_),
    .A2(_0989_),
    .B1(_1031_),
    .C1(_0813_),
    .Y(_1032_));
 sky130_fd_sc_hs__a21oi_4 _6039_ (.A1(_0814_),
    .A2(net92),
    .B1(_1032_),
    .Y(_1033_));
 sky130_fd_sc_hs__nor2_8 _6040_ (.A(_0109_),
    .B(_1033_),
    .Y(net268));
 sky130_fd_sc_hs__nand2_1 _6041_ (.A(_0814_),
    .B(net93),
    .Y(_1034_));
 sky130_fd_sc_hs__buf_4 _6042_ (.A(_0992_),
    .X(_1035_));
 sky130_fd_sc_hs__nand2b_1 _6043_ (.A_N(net165),
    .B(_1035_),
    .Y(_1036_));
 sky130_fd_sc_hs__buf_8 _6044_ (.A(_0090_),
    .X(_1037_));
 sky130_fd_sc_hs__o211ai_2 _6045_ (.A1(net203),
    .A2(_0993_),
    .B1(_1036_),
    .C1(_1037_),
    .Y(_1038_));
 sky130_fd_sc_hs__a21oi_4 _6046_ (.A1(_1034_),
    .A2(_1038_),
    .B1(_0109_),
    .Y(net269));
 sky130_fd_sc_hs__buf_4 _6047_ (.A(_0989_),
    .X(_1039_));
 sky130_fd_sc_hs__nand2_1 _6048_ (.A(net204),
    .B(_1039_),
    .Y(_1040_));
 sky130_fd_sc_hs__nand2_1 _6049_ (.A(net166),
    .B(_1013_),
    .Y(_1041_));
 sky130_fd_sc_hs__nor2_1 _6050_ (.A(_1029_),
    .B(net94),
    .Y(_1042_));
 sky130_fd_sc_hs__a311oi_4 _6051_ (.A1(_1023_),
    .A2(_1040_),
    .A3(_1041_),
    .B1(_1042_),
    .C1(_1019_),
    .Y(net270));
 sky130_fd_sc_hs__nand2_1 _6052_ (.A(net205),
    .B(_1039_),
    .Y(_1043_));
 sky130_fd_sc_hs__nand2_1 _6053_ (.A(net167),
    .B(_1013_),
    .Y(_1044_));
 sky130_fd_sc_hs__nor2_1 _6054_ (.A(_1029_),
    .B(net95),
    .Y(_1045_));
 sky130_fd_sc_hs__a311oi_4 _6055_ (.A1(_1023_),
    .A2(_1043_),
    .A3(_1044_),
    .B1(_1045_),
    .C1(_1019_),
    .Y(net271));
 sky130_fd_sc_hs__nand2_1 _6056_ (.A(net206),
    .B(_1039_),
    .Y(_1046_));
 sky130_fd_sc_hs__nand2_1 _6057_ (.A(net168),
    .B(_1013_),
    .Y(_1047_));
 sky130_fd_sc_hs__nor2_1 _6058_ (.A(_1029_),
    .B(net96),
    .Y(_1048_));
 sky130_fd_sc_hs__a311oi_4 _6059_ (.A1(_1023_),
    .A2(_1046_),
    .A3(_1047_),
    .B1(_1048_),
    .C1(_1019_),
    .Y(net272));
 sky130_fd_sc_hs__nand2_1 _6060_ (.A(net14),
    .B(_1039_),
    .Y(_1049_));
 sky130_fd_sc_hs__nand2_1 _6061_ (.A(net169),
    .B(_1013_),
    .Y(_1050_));
 sky130_fd_sc_hs__nor2_1 _6062_ (.A(_1029_),
    .B(net97),
    .Y(_1051_));
 sky130_fd_sc_hs__a311oi_4 _6063_ (.A1(_1023_),
    .A2(_1049_),
    .A3(_1050_),
    .B1(_1051_),
    .C1(_1019_),
    .Y(net273));
 sky130_fd_sc_hs__nand2_1 _6064_ (.A(net208),
    .B(_1039_),
    .Y(_1052_));
 sky130_fd_sc_hs__nand2_1 _6065_ (.A(net170),
    .B(_1013_),
    .Y(_1053_));
 sky130_fd_sc_hs__nor2_1 _6066_ (.A(_1029_),
    .B(net98),
    .Y(_1054_));
 sky130_fd_sc_hs__a311oi_4 _6067_ (.A1(_1023_),
    .A2(_1052_),
    .A3(_1053_),
    .B1(_1054_),
    .C1(_1019_),
    .Y(net274));
 sky130_fd_sc_hs__nand2_1 _6068_ (.A(net209),
    .B(_1039_),
    .Y(_1055_));
 sky130_fd_sc_hs__nand2_1 _6069_ (.A(net171),
    .B(_1035_),
    .Y(_1056_));
 sky130_fd_sc_hs__nor2_1 _6070_ (.A(_1029_),
    .B(net99),
    .Y(_1057_));
 sky130_fd_sc_hs__a311oi_4 _6071_ (.A1(_1023_),
    .A2(_1055_),
    .A3(_1056_),
    .B1(_1057_),
    .C1(_1019_),
    .Y(net275));
 sky130_fd_sc_hs__nand2_1 _6072_ (.A(_0814_),
    .B(net100),
    .Y(_1058_));
 sky130_fd_sc_hs__nand2b_1 _6073_ (.A_N(net172),
    .B(_0992_),
    .Y(_1059_));
 sky130_fd_sc_hs__o211ai_2 _6074_ (.A1(net210),
    .A2(_0993_),
    .B1(_1059_),
    .C1(_1037_),
    .Y(_1060_));
 sky130_fd_sc_hs__a21oi_4 _6075_ (.A1(_1058_),
    .A2(_1060_),
    .B1(_0109_),
    .Y(net276));
 sky130_fd_sc_hs__nand2_1 _6076_ (.A(net12),
    .B(_1039_),
    .Y(_1061_));
 sky130_fd_sc_hs__nand2_1 _6077_ (.A(net173),
    .B(_1035_),
    .Y(_1062_));
 sky130_fd_sc_hs__nor2_1 _6078_ (.A(_1029_),
    .B(net101),
    .Y(_1063_));
 sky130_fd_sc_hs__a311oi_4 _6079_ (.A1(_1023_),
    .A2(_1061_),
    .A3(_1062_),
    .B1(_1063_),
    .C1(_0600_),
    .Y(net277));
 sky130_fd_sc_hs__nand2_1 _6080_ (.A(net9),
    .B(_1039_),
    .Y(_1064_));
 sky130_fd_sc_hs__nand2_1 _6081_ (.A(net174),
    .B(_1035_),
    .Y(_1065_));
 sky130_fd_sc_hs__nor2_1 _6082_ (.A(_1029_),
    .B(net102),
    .Y(_1066_));
 sky130_fd_sc_hs__a311oi_4 _6083_ (.A1(_1023_),
    .A2(_1064_),
    .A3(_1065_),
    .B1(_1066_),
    .C1(_0600_),
    .Y(net278));
 sky130_fd_sc_hs__nand2_1 _6084_ (.A(net213),
    .B(_1039_),
    .Y(_1067_));
 sky130_fd_sc_hs__nand2_1 _6085_ (.A(net175),
    .B(_1035_),
    .Y(_1068_));
 sky130_fd_sc_hs__nor2_1 _6086_ (.A(_1029_),
    .B(net103),
    .Y(_1069_));
 sky130_fd_sc_hs__a311oi_4 _6087_ (.A1(_1037_),
    .A2(_1067_),
    .A3(_1068_),
    .B1(_1069_),
    .C1(_0600_),
    .Y(net279));
 sky130_fd_sc_hs__nand2_1 _6088_ (.A(_0814_),
    .B(net104),
    .Y(_1070_));
 sky130_fd_sc_hs__nand2b_1 _6089_ (.A_N(net176),
    .B(_0992_),
    .Y(_1071_));
 sky130_fd_sc_hs__o211ai_2 _6090_ (.A1(net214),
    .A2(_0993_),
    .B1(_1071_),
    .C1(_1037_),
    .Y(_1072_));
 sky130_fd_sc_hs__a21oi_4 _6091_ (.A1(_1070_),
    .A2(_1072_),
    .B1(_0109_),
    .Y(net280));
 sky130_fd_sc_hs__nand2_1 _6092_ (.A(_0814_),
    .B(net105),
    .Y(_1073_));
 sky130_fd_sc_hs__o211ai_4 _6093_ (.A1(_0523_),
    .A2(net215),
    .B1(_1037_),
    .C1(net177),
    .Y(_1074_));
 sky130_fd_sc_hs__a21oi_4 _6094_ (.A1(_1073_),
    .A2(_1074_),
    .B1(_0109_),
    .Y(net281));
 sky130_fd_sc_hs__nand2b_4 _6095_ (.A_N(net185),
    .B(net186),
    .Y(_1075_));
 sky130_fd_sc_hs__buf_8 _6096_ (.A(_1075_),
    .X(_1076_));
 sky130_fd_sc_hs__buf_8 _6097_ (.A(_1076_),
    .X(_1077_));
 sky130_fd_sc_hs__mux2i_4 _6098_ (.A0(_0435_),
    .A1(net191),
    .S(_0959_),
    .Y(_1078_));
 sky130_fd_sc_hs__buf_8 _6099_ (.A(_1076_),
    .X(_1079_));
 sky130_fd_sc_hs__a211oi_4 _6100_ (.A1(_0920_),
    .A2(_0977_),
    .B1(_1079_),
    .C1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[0] ),
    .Y(_1080_));
 sky130_fd_sc_hs__nand2_4 _6101_ (.A(_0105_),
    .B(_0386_),
    .Y(_1081_));
 sky130_fd_sc_hs__buf_8 _6102_ (.A(_1081_),
    .X(_1082_));
 sky130_fd_sc_hs__a211oi_4 _6103_ (.A1(_1077_),
    .A2(_1078_),
    .B1(_1080_),
    .C1(_1082_),
    .Y(_1083_));
 sky130_fd_sc_hs__nand2b_4 _6104_ (.A_N(net80),
    .B(_0104_),
    .Y(_1084_));
 sky130_fd_sc_hs__buf_8 _6105_ (.A(_1084_),
    .X(_1085_));
 sky130_fd_sc_hs__buf_8 _6106_ (.A(_1085_),
    .X(_1086_));
 sky130_fd_sc_hs__nor2_4 _6107_ (.A(_0081_),
    .B(\genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0] ),
    .Y(_1087_));
 sky130_fd_sc_hs__nand2_8 _6108_ (.A(_0083_),
    .B(_1087_),
    .Y(_1088_));
 sky130_fd_sc_hs__buf_8 _6109_ (.A(_1088_),
    .X(_1089_));
 sky130_fd_sc_hs__mux2i_4 _6110_ (.A0(_0435_),
    .A1(_3701_),
    .S(_1089_),
    .Y(_1090_));
 sky130_fd_sc_hs__mux4_1 _6111_ (.A0(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[31] ),
    .A1(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[30] ),
    .A2(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[29] ),
    .A3(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[28] ),
    .S0(_0590_),
    .S1(_0823_),
    .X(_1091_));
 sky130_fd_sc_hs__mux4_1 _6112_ (.A0(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[27] ),
    .A1(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[26] ),
    .A2(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[25] ),
    .A3(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[24] ),
    .S0(_0590_),
    .S1(_0823_),
    .X(_1092_));
 sky130_fd_sc_hs__mux4_1 _6113_ (.A0(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[23] ),
    .A1(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[22] ),
    .A2(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[21] ),
    .A3(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[20] ),
    .S0(_0590_),
    .S1(_0823_),
    .X(_1093_));
 sky130_fd_sc_hs__mux4_1 _6114_ (.A0(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[19] ),
    .A1(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[18] ),
    .A2(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[17] ),
    .A3(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[16] ),
    .S0(_0589_),
    .S1(_0823_),
    .X(_1094_));
 sky130_fd_sc_hs__xnor2_4 _6115_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .B(_3706_),
    .Y(_1095_));
 sky130_fd_sc_hs__mux4_4 _6116_ (.A0(_1091_),
    .A1(_1092_),
    .A2(_1093_),
    .A3(_1094_),
    .S0(_1095_),
    .S1(_0828_),
    .X(_1096_));
 sky130_fd_sc_hs__mux4_1 _6117_ (.A0(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[15] ),
    .A1(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[14] ),
    .A2(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[13] ),
    .A3(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[12] ),
    .S0(_0590_),
    .S1(_0823_),
    .X(_1097_));
 sky130_fd_sc_hs__mux4_1 _6118_ (.A0(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[11] ),
    .A1(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[10] ),
    .A2(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[9] ),
    .A3(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[8] ),
    .S0(_0590_),
    .S1(_0823_),
    .X(_1098_));
 sky130_fd_sc_hs__mux4_1 _6119_ (.A0(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[7] ),
    .A1(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[6] ),
    .A2(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[5] ),
    .A3(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[4] ),
    .S0(_0590_),
    .S1(_0823_),
    .X(_1099_));
 sky130_fd_sc_hs__mux4_1 _6120_ (.A0(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[3] ),
    .A1(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[2] ),
    .A2(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[1] ),
    .A3(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[0] ),
    .S0(_0589_),
    .S1(_0823_),
    .X(_1100_));
 sky130_fd_sc_hs__mux4_2 _6121_ (.A0(_1097_),
    .A1(_1098_),
    .A2(_1099_),
    .A3(_1100_),
    .S0(_1095_),
    .S1(_0828_),
    .X(_1101_));
 sky130_fd_sc_hs__xnor2_4 _6122_ (.A(_0096_),
    .B(_0829_),
    .Y(_1102_));
 sky130_fd_sc_hs__mux2i_4 _6123_ (.A0(_1096_),
    .A1(_1101_),
    .S(_1102_),
    .Y(_1103_));
 sky130_fd_sc_hs__nor3_2 _6124_ (.A(_0513_),
    .B(_0992_),
    .C(_1075_),
    .Y(_1104_));
 sky130_fd_sc_hs__a21oi_4 _6125_ (.A1(_0513_),
    .A2(_0992_),
    .B1(_1104_),
    .Y(_1105_));
 sky130_fd_sc_hs__o22ai_4 _6126_ (.A1(_0841_),
    .A2(_0818_),
    .B1(_1105_),
    .B2(\genblk3.gen_multdiv_fast.multdiv_i.div_by_zero_q ),
    .Y(_1106_));
 sky130_fd_sc_hs__clkbuf_8 _6127_ (.A(_1106_),
    .X(_1107_));
 sky130_fd_sc_hs__mux2i_1 _6128_ (.A0(_0435_),
    .A1(net191),
    .S(_1107_),
    .Y(_1108_));
 sky130_fd_sc_hs__buf_8 _6129_ (.A(_0381_),
    .X(_1109_));
 sky130_fd_sc_hs__or4_4 _6130_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.md_state_q[2] ),
    .B(_0378_),
    .C(\genblk3.gen_multdiv_fast.multdiv_i.md_state_q[0] ),
    .D(_0393_),
    .X(_1110_));
 sky130_fd_sc_hs__nand2_8 _6131_ (.A(_0819_),
    .B(_1110_),
    .Y(_1111_));
 sky130_fd_sc_hs__a221oi_4 _6132_ (.A1(net121),
    .A2(_0122_),
    .B1(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[31] ),
    .B2(_0090_),
    .C1(_1111_),
    .Y(_1112_));
 sky130_fd_sc_hs__o221a_1 _6133_ (.A1(_0391_),
    .A2(_1103_),
    .B1(_1108_),
    .B2(_1109_),
    .C1(_1112_),
    .X(_1113_));
 sky130_fd_sc_hs__clkbuf_8 _6134_ (.A(_1110_),
    .X(_1114_));
 sky130_fd_sc_hs__buf_4 _6135_ (.A(_1114_),
    .X(_1115_));
 sky130_fd_sc_hs__clkbuf_8 _6136_ (.A(_0105_),
    .X(_1116_));
 sky130_fd_sc_hs__o21ai_1 _6137_ (.A1(_0435_),
    .A2(_1115_),
    .B1(_1116_),
    .Y(_1117_));
 sky130_fd_sc_hs__o22ai_1 _6138_ (.A1(_1086_),
    .A2(_1090_),
    .B1(_1113_),
    .B2(_1117_),
    .Y(_1118_));
 sky130_fd_sc_hs__or2_1 _6139_ (.A(_1083_),
    .B(_1118_),
    .X(net282));
 sky130_fd_sc_hs__nor2b_4 _6140_ (.A(_0105_),
    .B_N(_0104_),
    .Y(_1119_));
 sky130_fd_sc_hs__mux2_2 _6141_ (.A0(_0447_),
    .A1(_3716_),
    .S(_1088_),
    .X(_1120_));
 sky130_fd_sc_hs__nand2_8 _6142_ (.A(_1119_),
    .B(_1120_),
    .Y(_1121_));
 sky130_fd_sc_hs__clkbuf_8 _6143_ (.A(_1114_),
    .X(_1122_));
 sky130_fd_sc_hs__buf_4 _6144_ (.A(_0105_),
    .X(_1123_));
 sky130_fd_sc_hs__o21ai_2 _6145_ (.A1(_0447_),
    .A2(_1122_),
    .B1(_1123_),
    .Y(_1124_));
 sky130_fd_sc_hs__buf_8 _6146_ (.A(_0818_),
    .X(_1125_));
 sky130_fd_sc_hs__buf_8 _6147_ (.A(_1125_),
    .X(_1126_));
 sky130_fd_sc_hs__clkbuf_16 _6148_ (.A(_0958_),
    .X(_1127_));
 sky130_fd_sc_hs__mux2_1 _6149_ (.A0(_0447_),
    .A1(net202),
    .S(_1127_),
    .X(_1128_));
 sky130_fd_sc_hs__buf_8 _6150_ (.A(_1076_),
    .X(_1129_));
 sky130_fd_sc_hs__a211o_1 _6151_ (.A1(_0100_),
    .A2(_0959_),
    .B1(_1129_),
    .C1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[1] ),
    .X(_1130_));
 sky130_fd_sc_hs__o211ai_2 _6152_ (.A1(_1126_),
    .A2(_1128_),
    .B1(_1130_),
    .C1(_0386_),
    .Y(_1131_));
 sky130_fd_sc_hs__buf_8 _6153_ (.A(_1111_),
    .X(_1132_));
 sky130_fd_sc_hs__a21oi_4 _6154_ (.A1(net132),
    .A2(_0123_),
    .B1(_1132_),
    .Y(_1133_));
 sky130_fd_sc_hs__buf_8 _6155_ (.A(_1106_),
    .X(_1134_));
 sky130_fd_sc_hs__nand2_1 _6156_ (.A(_0306_),
    .B(_1134_),
    .Y(_1135_));
 sky130_fd_sc_hs__o211ai_1 _6157_ (.A1(_0447_),
    .A2(_1134_),
    .B1(_1135_),
    .C1(_0430_),
    .Y(_1136_));
 sky130_fd_sc_hs__o2111a_1 _6158_ (.A1(_0433_),
    .A2(_1078_),
    .B1(_1121_),
    .C1(_1133_),
    .D1(_1136_),
    .X(_1137_));
 sky130_fd_sc_hs__a22oi_4 _6159_ (.A1(_1121_),
    .A2(_1124_),
    .B1(_1131_),
    .B2(_1137_),
    .Y(net283));
 sky130_fd_sc_hs__nor2_1 _6160_ (.A(_0314_),
    .B(_0932_),
    .Y(_1138_));
 sky130_fd_sc_hs__a21oi_4 _6161_ (.A1(_0450_),
    .A2(_0932_),
    .B1(_1138_),
    .Y(_1139_));
 sky130_fd_sc_hs__a211oi_4 _6162_ (.A1(_0938_),
    .A2(_0977_),
    .B1(_1076_),
    .C1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[2] ),
    .Y(_1140_));
 sky130_fd_sc_hs__a211oi_4 _6163_ (.A1(_1129_),
    .A2(_1139_),
    .B1(_1140_),
    .C1(_1082_),
    .Y(_1141_));
 sky130_fd_sc_hs__and2_4 _6164_ (.A(_0083_),
    .B(_1087_),
    .X(_1142_));
 sky130_fd_sc_hs__buf_4 _6165_ (.A(_1142_),
    .X(_1143_));
 sky130_fd_sc_hs__clkbuf_8 _6166_ (.A(_1143_),
    .X(_1144_));
 sky130_fd_sc_hs__nand2_1 _6167_ (.A(_0450_),
    .B(_1144_),
    .Y(_1145_));
 sky130_fd_sc_hs__clkbuf_8 _6168_ (.A(_1088_),
    .X(_1146_));
 sky130_fd_sc_hs__buf_8 _6169_ (.A(_1146_),
    .X(_1147_));
 sky130_fd_sc_hs__nand2_1 _6170_ (.A(_3718_),
    .B(_1147_),
    .Y(_1148_));
 sky130_fd_sc_hs__a21oi_1 _6171_ (.A1(_1145_),
    .A2(_1148_),
    .B1(_1086_),
    .Y(_1149_));
 sky130_fd_sc_hs__nand2_1 _6172_ (.A(_0103_),
    .B(_1128_),
    .Y(_1150_));
 sky130_fd_sc_hs__buf_8 _6173_ (.A(_1106_),
    .X(_1151_));
 sky130_fd_sc_hs__mux2i_1 _6174_ (.A0(_0450_),
    .A1(net213),
    .S(_1151_),
    .Y(_1152_));
 sky130_fd_sc_hs__buf_8 _6175_ (.A(_0122_),
    .X(_1153_));
 sky130_fd_sc_hs__buf_8 _6176_ (.A(_1111_),
    .X(_1154_));
 sky130_fd_sc_hs__a21oi_1 _6177_ (.A1(net143),
    .A2(_1153_),
    .B1(_1154_),
    .Y(_1155_));
 sky130_fd_sc_hs__o21a_1 _6178_ (.A1(_1109_),
    .A2(_1152_),
    .B1(_1155_),
    .X(_1156_));
 sky130_fd_sc_hs__o21ai_1 _6179_ (.A1(_0450_),
    .A2(_1115_),
    .B1(_1116_),
    .Y(_1157_));
 sky130_fd_sc_hs__a21oi_1 _6180_ (.A1(_1150_),
    .A2(_1156_),
    .B1(_1157_),
    .Y(_1158_));
 sky130_fd_sc_hs__or3_2 _6181_ (.A(_1141_),
    .B(_1149_),
    .C(_1158_),
    .X(net284));
 sky130_fd_sc_hs__nand2_1 _6182_ (.A(_0572_),
    .B(_1142_),
    .Y(_1159_));
 sky130_fd_sc_hs__nand2_1 _6183_ (.A(_3726_),
    .B(_1088_),
    .Y(_1160_));
 sky130_fd_sc_hs__a21oi_4 _6184_ (.A1(_1159_),
    .A2(_1160_),
    .B1(_1085_),
    .Y(_1161_));
 sky130_fd_sc_hs__o21a_1 _6185_ (.A1(_0572_),
    .A2(_1122_),
    .B1(_1123_),
    .X(_1162_));
 sky130_fd_sc_hs__mux2i_1 _6186_ (.A0(_0572_),
    .A1(net216),
    .S(_1134_),
    .Y(_1163_));
 sky130_fd_sc_hs__clkbuf_16 _6187_ (.A(_0122_),
    .X(_1164_));
 sky130_fd_sc_hs__a211oi_4 _6188_ (.A1(net146),
    .A2(_1164_),
    .B1(_1154_),
    .C1(_1161_),
    .Y(_1165_));
 sky130_fd_sc_hs__o221a_1 _6189_ (.A1(_0433_),
    .A2(_1139_),
    .B1(_1163_),
    .B2(_0810_),
    .C1(_1165_),
    .X(_1166_));
 sky130_fd_sc_hs__mux2i_4 _6190_ (.A0(_0572_),
    .A1(net216),
    .S(_1127_),
    .Y(_1167_));
 sky130_fd_sc_hs__a311oi_4 _6191_ (.A1(_0941_),
    .A2(_0099_),
    .A3(_0959_),
    .B1(_1079_),
    .C1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[3] ),
    .Y(_1168_));
 sky130_fd_sc_hs__a21oi_1 _6192_ (.A1(_1077_),
    .A2(_1167_),
    .B1(_1168_),
    .Y(_1169_));
 sky130_fd_sc_hs__nand2_1 _6193_ (.A(_0386_),
    .B(_1169_),
    .Y(_1170_));
 sky130_fd_sc_hs__a2bb2oi_4 _6194_ (.A1_N(_1161_),
    .A2_N(_1162_),
    .B1(_1166_),
    .B2(_1170_),
    .Y(net285));
 sky130_fd_sc_hs__a211oi_4 _6195_ (.A1(_0920_),
    .A2(_0984_),
    .B1(_1077_),
    .C1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[4] ),
    .Y(_1171_));
 sky130_fd_sc_hs__mux2_1 _6196_ (.A0(_0573_),
    .A1(net217),
    .S(_1127_),
    .X(_1172_));
 sky130_fd_sc_hs__nor2_2 _6197_ (.A(_1126_),
    .B(_1172_),
    .Y(_1173_));
 sky130_fd_sc_hs__mux2i_1 _6198_ (.A0(_0573_),
    .A1(net217),
    .S(_1151_),
    .Y(_1174_));
 sky130_fd_sc_hs__a21oi_4 _6199_ (.A1(net147),
    .A2(_0123_),
    .B1(_1132_),
    .Y(_1175_));
 sky130_fd_sc_hs__o221ai_1 _6200_ (.A1(_0433_),
    .A2(_1167_),
    .B1(_1174_),
    .B2(_0810_),
    .C1(_1175_),
    .Y(_1176_));
 sky130_fd_sc_hs__o21a_1 _6201_ (.A1(_0573_),
    .A2(_1115_),
    .B1(_1116_),
    .X(_1177_));
 sky130_fd_sc_hs__buf_8 _6202_ (.A(_1143_),
    .X(_1178_));
 sky130_fd_sc_hs__nand2_1 _6203_ (.A(_0573_),
    .B(_1178_),
    .Y(_1179_));
 sky130_fd_sc_hs__nand2_1 _6204_ (.A(_3730_),
    .B(_1147_),
    .Y(_1180_));
 sky130_fd_sc_hs__a21oi_2 _6205_ (.A1(_1179_),
    .A2(_1180_),
    .B1(_1086_),
    .Y(_1181_));
 sky130_fd_sc_hs__a21oi_2 _6206_ (.A1(_1176_),
    .A2(_1177_),
    .B1(_1181_),
    .Y(_1182_));
 sky130_fd_sc_hs__o31ai_4 _6207_ (.A1(_1082_),
    .A2(_1171_),
    .A3(_1173_),
    .B1(_1182_),
    .Y(net286));
 sky130_fd_sc_hs__nor2_1 _6208_ (.A(_0317_),
    .B(_0932_),
    .Y(_1183_));
 sky130_fd_sc_hs__a21oi_4 _6209_ (.A1(_0574_),
    .A2(_0932_),
    .B1(_1183_),
    .Y(_1184_));
 sky130_fd_sc_hs__a211oi_4 _6210_ (.A1(_0095_),
    .A2(_0984_),
    .B1(_1076_),
    .C1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[5] ),
    .Y(_1185_));
 sky130_fd_sc_hs__a211oi_4 _6211_ (.A1(_1129_),
    .A2(_1184_),
    .B1(_1185_),
    .C1(_1082_),
    .Y(_1186_));
 sky130_fd_sc_hs__nand2_1 _6212_ (.A(_0574_),
    .B(_1144_),
    .Y(_1187_));
 sky130_fd_sc_hs__nand2_1 _6213_ (.A(_3739_),
    .B(_1147_),
    .Y(_1188_));
 sky130_fd_sc_hs__a21oi_1 _6214_ (.A1(_1187_),
    .A2(_1188_),
    .B1(_1086_),
    .Y(_1189_));
 sky130_fd_sc_hs__nand2_1 _6215_ (.A(_0103_),
    .B(_1172_),
    .Y(_1190_));
 sky130_fd_sc_hs__a2bb2oi_4 _6216_ (.A1_N(\genblk3.gen_multdiv_fast.multdiv_i.div_by_zero_q ),
    .A2_N(_1105_),
    .B1(_1075_),
    .B2(_0835_),
    .Y(_1191_));
 sky130_fd_sc_hs__buf_8 _6217_ (.A(_1191_),
    .X(_1192_));
 sky130_fd_sc_hs__nor2_1 _6218_ (.A(_0317_),
    .B(_1191_),
    .Y(_1193_));
 sky130_fd_sc_hs__a21oi_1 _6219_ (.A1(_0574_),
    .A2(_1192_),
    .B1(_1193_),
    .Y(_1194_));
 sky130_fd_sc_hs__a21oi_1 _6220_ (.A1(net148),
    .A2(_1153_),
    .B1(_1154_),
    .Y(_1195_));
 sky130_fd_sc_hs__o21a_1 _6221_ (.A1(_1109_),
    .A2(_1194_),
    .B1(_1195_),
    .X(_1196_));
 sky130_fd_sc_hs__o21ai_1 _6222_ (.A1(_0574_),
    .A2(_1115_),
    .B1(_1116_),
    .Y(_1197_));
 sky130_fd_sc_hs__a21oi_1 _6223_ (.A1(_1190_),
    .A2(_1196_),
    .B1(_1197_),
    .Y(_1198_));
 sky130_fd_sc_hs__or3_4 _6224_ (.A(_1186_),
    .B(_1189_),
    .C(_1198_),
    .X(net287));
 sky130_fd_sc_hs__nand2_1 _6225_ (.A(net216),
    .B(_1039_),
    .Y(_1199_));
 sky130_fd_sc_hs__nand2_1 _6226_ (.A(net178),
    .B(_1035_),
    .Y(_1200_));
 sky130_fd_sc_hs__nor2_1 _6227_ (.A(_0090_),
    .B(net106),
    .Y(_1201_));
 sky130_fd_sc_hs__a311oi_4 _6228_ (.A1(_1037_),
    .A2(_1199_),
    .A3(_1200_),
    .B1(_1201_),
    .C1(_0600_),
    .Y(net288));
 sky130_fd_sc_hs__nand2_1 _6229_ (.A(_0575_),
    .B(_1142_),
    .Y(_1202_));
 sky130_fd_sc_hs__nand2_1 _6230_ (.A(_3749_),
    .B(_1088_),
    .Y(_1203_));
 sky130_fd_sc_hs__a21oi_4 _6231_ (.A1(_1202_),
    .A2(_1203_),
    .B1(_1085_),
    .Y(_1204_));
 sky130_fd_sc_hs__o21a_1 _6232_ (.A1(_0575_),
    .A2(_1122_),
    .B1(_1123_),
    .X(_1205_));
 sky130_fd_sc_hs__mux2i_1 _6233_ (.A0(_0575_),
    .A1(net219),
    .S(_1134_),
    .Y(_1206_));
 sky130_fd_sc_hs__a211oi_4 _6234_ (.A1(net149),
    .A2(_1164_),
    .B1(_1154_),
    .C1(_1204_),
    .Y(_1207_));
 sky130_fd_sc_hs__o221a_2 _6235_ (.A1(_0433_),
    .A2(_1184_),
    .B1(_1206_),
    .B2(_0810_),
    .C1(_1207_),
    .X(_1208_));
 sky130_fd_sc_hs__a211oi_4 _6236_ (.A1(_0938_),
    .A2(_0984_),
    .B1(_1079_),
    .C1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[6] ),
    .Y(_1209_));
 sky130_fd_sc_hs__clkbuf_8 _6237_ (.A(_0818_),
    .X(_1210_));
 sky130_fd_sc_hs__clkbuf_16 _6238_ (.A(_0958_),
    .X(_1211_));
 sky130_fd_sc_hs__mux2_1 _6239_ (.A0(_0575_),
    .A1(net219),
    .S(_1211_),
    .X(_1212_));
 sky130_fd_sc_hs__nor2_1 _6240_ (.A(_1210_),
    .B(_1212_),
    .Y(_1213_));
 sky130_fd_sc_hs__or3_1 _6241_ (.A(_0392_),
    .B(_1209_),
    .C(_1213_),
    .X(_1214_));
 sky130_fd_sc_hs__a2bb2oi_4 _6242_ (.A1_N(_1204_),
    .A2_N(_1205_),
    .B1(_1208_),
    .B2(_1214_),
    .Y(net289));
 sky130_fd_sc_hs__nand2_1 _6243_ (.A(_0576_),
    .B(_1142_),
    .Y(_1215_));
 sky130_fd_sc_hs__nand2_1 _6244_ (.A(_2347_),
    .B(_1088_),
    .Y(_1216_));
 sky130_fd_sc_hs__a21oi_4 _6245_ (.A1(_1215_),
    .A2(_1216_),
    .B1(_1085_),
    .Y(_1217_));
 sky130_fd_sc_hs__o21a_1 _6246_ (.A1(_0576_),
    .A2(_1122_),
    .B1(_1123_),
    .X(_1218_));
 sky130_fd_sc_hs__mux2i_4 _6247_ (.A0(_0576_),
    .A1(net220),
    .S(_1134_),
    .Y(_1219_));
 sky130_fd_sc_hs__a211oi_4 _6248_ (.A1(net150),
    .A2(_1164_),
    .B1(_1154_),
    .C1(_1217_),
    .Y(_1220_));
 sky130_fd_sc_hs__o21ai_4 _6249_ (.A1(_0810_),
    .A2(_1219_),
    .B1(_1220_),
    .Y(_1221_));
 sky130_fd_sc_hs__a21oi_1 _6250_ (.A1(_0103_),
    .A2(_1212_),
    .B1(_1221_),
    .Y(_1222_));
 sky130_fd_sc_hs__a211oi_4 _6251_ (.A1(_0941_),
    .A2(_0984_),
    .B1(_1079_),
    .C1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[7] ),
    .Y(_1223_));
 sky130_fd_sc_hs__mux2_4 _6252_ (.A0(_0576_),
    .A1(net220),
    .S(_1127_),
    .X(_1224_));
 sky130_fd_sc_hs__nor2_1 _6253_ (.A(_1210_),
    .B(_1224_),
    .Y(_1225_));
 sky130_fd_sc_hs__or3_1 _6254_ (.A(_0392_),
    .B(_1223_),
    .C(_1225_),
    .X(_1226_));
 sky130_fd_sc_hs__a2bb2oi_2 _6255_ (.A1_N(_1217_),
    .A2_N(_1218_),
    .B1(_1222_),
    .B2(_1226_),
    .Y(net290));
 sky130_fd_sc_hs__mux2_1 _6256_ (.A0(_0577_),
    .A1(net221),
    .S(_1151_),
    .X(_1227_));
 sky130_fd_sc_hs__nor2_2 _6257_ (.A(net151),
    .B(_1125_),
    .Y(_1228_));
 sky130_fd_sc_hs__nor2_8 _6258_ (.A(_0392_),
    .B(_1075_),
    .Y(_1229_));
 sky130_fd_sc_hs__a21oi_4 _6259_ (.A1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[8] ),
    .A2(_1229_),
    .B1(_1164_),
    .Y(_1230_));
 sky130_fd_sc_hs__buf_8 _6260_ (.A(_1114_),
    .X(_1231_));
 sky130_fd_sc_hs__xnor2_4 _6261_ (.A(_3766_),
    .B(_2346_),
    .Y(_1232_));
 sky130_fd_sc_hs__nand2_1 _6262_ (.A(_1146_),
    .B(_1232_),
    .Y(_1233_));
 sky130_fd_sc_hs__o211ai_4 _6263_ (.A1(_0577_),
    .A2(_1146_),
    .B1(_1233_),
    .C1(_1119_),
    .Y(_1234_));
 sky130_fd_sc_hs__o211ai_4 _6264_ (.A1(_1228_),
    .A2(_1230_),
    .B1(_1231_),
    .C1(_1234_),
    .Y(_1235_));
 sky130_fd_sc_hs__a221oi_4 _6265_ (.A1(_0103_),
    .A2(_1224_),
    .B1(_1227_),
    .B2(_0430_),
    .C1(_1235_),
    .Y(_1236_));
 sky130_fd_sc_hs__mux2i_4 _6266_ (.A0(_0577_),
    .A1(net221),
    .S(_1211_),
    .Y(_1237_));
 sky130_fd_sc_hs__nor2_1 _6267_ (.A(_1210_),
    .B(_1237_),
    .Y(_1238_));
 sky130_fd_sc_hs__and3_1 _6268_ (.A(_0920_),
    .B(_1125_),
    .C(_0937_),
    .X(_1239_));
 sky130_fd_sc_hs__o21ai_1 _6269_ (.A1(_1238_),
    .A2(_1239_),
    .B1(_0386_),
    .Y(_1240_));
 sky130_fd_sc_hs__clkbuf_8 _6270_ (.A(_0105_),
    .X(_1241_));
 sky130_fd_sc_hs__buf_8 _6271_ (.A(_1241_),
    .X(_1242_));
 sky130_fd_sc_hs__o21ai_1 _6272_ (.A1(_0577_),
    .A2(_1122_),
    .B1(_1242_),
    .Y(_1243_));
 sky130_fd_sc_hs__a22oi_4 _6273_ (.A1(_1236_),
    .A2(_1240_),
    .B1(_1243_),
    .B2(_1234_),
    .Y(net291));
 sky130_fd_sc_hs__a21oi_1 _6274_ (.A1(_0095_),
    .A2(_0937_),
    .B1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[9] ),
    .Y(_1244_));
 sky130_fd_sc_hs__mux2_1 _6275_ (.A0(_0578_),
    .A1(net222),
    .S(_0958_),
    .X(_1245_));
 sky130_fd_sc_hs__o21ai_4 _6276_ (.A1(_0566_),
    .A2(_1114_),
    .B1(_0105_),
    .Y(_1246_));
 sky130_fd_sc_hs__nor2_8 _6277_ (.A(_0392_),
    .B(_1246_),
    .Y(_1247_));
 sky130_fd_sc_hs__o21ai_1 _6278_ (.A1(_1125_),
    .A2(_1245_),
    .B1(_1247_),
    .Y(_1248_));
 sky130_fd_sc_hs__a21oi_1 _6279_ (.A1(_1126_),
    .A2(_1244_),
    .B1(_1248_),
    .Y(_1249_));
 sky130_fd_sc_hs__nand2_1 _6280_ (.A(_0578_),
    .B(_1144_),
    .Y(_1250_));
 sky130_fd_sc_hs__a21o_1 _6281_ (.A1(_3756_),
    .A2(_2343_),
    .B1(_3755_),
    .X(_1251_));
 sky130_fd_sc_hs__a21oi_4 _6282_ (.A1(_3766_),
    .A2(_1251_),
    .B1(_3765_),
    .Y(_1252_));
 sky130_fd_sc_hs__xnor2_4 _6283_ (.A(_3777_),
    .B(_1252_),
    .Y(_1253_));
 sky130_fd_sc_hs__nand2_4 _6284_ (.A(_1089_),
    .B(_1253_),
    .Y(_1254_));
 sky130_fd_sc_hs__a21oi_4 _6285_ (.A1(_1250_),
    .A2(_1254_),
    .B1(_1086_),
    .Y(_1255_));
 sky130_fd_sc_hs__nand2_1 _6286_ (.A(_0299_),
    .B(_1107_),
    .Y(_1256_));
 sky130_fd_sc_hs__o211ai_1 _6287_ (.A1(_0578_),
    .A2(_1151_),
    .B1(_1256_),
    .C1(_0378_),
    .Y(_1257_));
 sky130_fd_sc_hs__a21oi_4 _6288_ (.A1(net152),
    .A2(_1153_),
    .B1(_1111_),
    .Y(_1258_));
 sky130_fd_sc_hs__o211ai_2 _6289_ (.A1(_0391_),
    .A2(_1237_),
    .B1(_1257_),
    .C1(_1258_),
    .Y(_1259_));
 sky130_fd_sc_hs__o211a_1 _6290_ (.A1(_0578_),
    .A2(_1231_),
    .B1(_1259_),
    .C1(_1123_),
    .X(_1260_));
 sky130_fd_sc_hs__or3_1 _6291_ (.A(_1249_),
    .B(_1255_),
    .C(_1260_),
    .X(net292));
 sky130_fd_sc_hs__a211oi_4 _6292_ (.A1(_0938_),
    .A2(_0937_),
    .B1(_1077_),
    .C1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[10] ),
    .Y(_1261_));
 sky130_fd_sc_hs__mux2_2 _6293_ (.A0(_0580_),
    .A1(net192),
    .S(_1127_),
    .X(_1262_));
 sky130_fd_sc_hs__o21ai_1 _6294_ (.A1(_1126_),
    .A2(_1262_),
    .B1(_1247_),
    .Y(_1263_));
 sky130_fd_sc_hs__clkbuf_8 _6295_ (.A(_0102_),
    .X(_1264_));
 sky130_fd_sc_hs__nor2_2 _6296_ (.A(_0580_),
    .B(_1151_),
    .Y(_1265_));
 sky130_fd_sc_hs__nor2_2 _6297_ (.A(net192),
    .B(_1192_),
    .Y(_1266_));
 sky130_fd_sc_hs__a21oi_2 _6298_ (.A1(net122),
    .A2(_1153_),
    .B1(_1111_),
    .Y(_1267_));
 sky130_fd_sc_hs__o31ai_4 _6299_ (.A1(_1109_),
    .A2(_1265_),
    .A3(_1266_),
    .B1(_1267_),
    .Y(_1268_));
 sky130_fd_sc_hs__a21oi_1 _6300_ (.A1(_1264_),
    .A2(_1245_),
    .B1(_1268_),
    .Y(_1269_));
 sky130_fd_sc_hs__o21ai_1 _6301_ (.A1(_0580_),
    .A2(_1115_),
    .B1(_1116_),
    .Y(_1270_));
 sky130_fd_sc_hs__nand2_1 _6302_ (.A(_0580_),
    .B(_1144_),
    .Y(_1271_));
 sky130_fd_sc_hs__a21o_1 _6303_ (.A1(_3766_),
    .A2(_2346_),
    .B1(_3765_),
    .X(_1272_));
 sky130_fd_sc_hs__a21oi_4 _6304_ (.A1(_3777_),
    .A2(_1272_),
    .B1(_3776_),
    .Y(_1273_));
 sky130_fd_sc_hs__xnor2_4 _6305_ (.A(_3786_),
    .B(_1273_),
    .Y(_1274_));
 sky130_fd_sc_hs__nand2_1 _6306_ (.A(_1146_),
    .B(_1274_),
    .Y(_1275_));
 sky130_fd_sc_hs__a21oi_4 _6307_ (.A1(_1271_),
    .A2(_1275_),
    .B1(_1085_),
    .Y(_1276_));
 sky130_fd_sc_hs__o21bai_1 _6308_ (.A1(_1269_),
    .A2(_1270_),
    .B1_N(_1276_),
    .Y(_1277_));
 sky130_fd_sc_hs__o21bai_2 _6309_ (.A1(_1261_),
    .A2(_1263_),
    .B1_N(_1277_),
    .Y(net293));
 sky130_fd_sc_hs__nand2_1 _6310_ (.A(_0581_),
    .B(_1143_),
    .Y(_1278_));
 sky130_fd_sc_hs__inv_1 _6311_ (.A(_3777_),
    .Y(_1279_));
 sky130_fd_sc_hs__o21bai_4 _6312_ (.A1(_1279_),
    .A2(_1252_),
    .B1_N(_3776_),
    .Y(_1280_));
 sky130_fd_sc_hs__a21oi_4 _6313_ (.A1(_3786_),
    .A2(_1280_),
    .B1(_3785_),
    .Y(_1281_));
 sky130_fd_sc_hs__xnor2_4 _6314_ (.A(_3792_),
    .B(_1281_),
    .Y(_1282_));
 sky130_fd_sc_hs__nand2_1 _6315_ (.A(_1146_),
    .B(_1282_),
    .Y(_1283_));
 sky130_fd_sc_hs__a21oi_4 _6316_ (.A1(_1278_),
    .A2(_1283_),
    .B1(_1085_),
    .Y(_1284_));
 sky130_fd_sc_hs__o21a_1 _6317_ (.A1(_0581_),
    .A2(_1122_),
    .B1(_1123_),
    .X(_1285_));
 sky130_fd_sc_hs__mux2i_4 _6318_ (.A0(_0581_),
    .A1(net365),
    .S(_1151_),
    .Y(_1286_));
 sky130_fd_sc_hs__a21oi_4 _6319_ (.A1(net123),
    .A2(_1164_),
    .B1(_1132_),
    .Y(_1287_));
 sky130_fd_sc_hs__o21ai_4 _6320_ (.A1(_0810_),
    .A2(_1286_),
    .B1(_1287_),
    .Y(_1288_));
 sky130_fd_sc_hs__a211oi_4 _6321_ (.A1(_0103_),
    .A2(_1262_),
    .B1(_1284_),
    .C1(_1288_),
    .Y(_1289_));
 sky130_fd_sc_hs__mux2i_4 _6322_ (.A0(_0581_),
    .A1(net365),
    .S(_0959_),
    .Y(_1290_));
 sky130_fd_sc_hs__a211oi_4 _6323_ (.A1(_0941_),
    .A2(_0937_),
    .B1(_1079_),
    .C1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[11] ),
    .Y(_1291_));
 sky130_fd_sc_hs__a211o_1 _6324_ (.A1(_1077_),
    .A2(_1290_),
    .B1(_1291_),
    .C1(_0392_),
    .X(_1292_));
 sky130_fd_sc_hs__a2bb2oi_4 _6325_ (.A1_N(_1284_),
    .A2_N(_1285_),
    .B1(_1289_),
    .B2(_1292_),
    .Y(net294));
 sky130_fd_sc_hs__mux2i_4 _6326_ (.A0(_0582_),
    .A1(net194),
    .S(_1211_),
    .Y(_1293_));
 sky130_fd_sc_hs__a211oi_4 _6327_ (.A1(_0920_),
    .A2(_0945_),
    .B1(_1076_),
    .C1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[12] ),
    .Y(_1294_));
 sky130_fd_sc_hs__a211oi_4 _6328_ (.A1(_1079_),
    .A2(_1293_),
    .B1(_1294_),
    .C1(_0392_),
    .Y(_1295_));
 sky130_fd_sc_hs__mux2i_4 _6329_ (.A0(_0582_),
    .A1(net194),
    .S(_1151_),
    .Y(_1296_));
 sky130_fd_sc_hs__nand2_1 _6330_ (.A(_0582_),
    .B(_1142_),
    .Y(_1297_));
 sky130_fd_sc_hs__inv_2 _6331_ (.A(_3801_),
    .Y(_1298_));
 sky130_fd_sc_hs__inv_2 _6332_ (.A(_3792_),
    .Y(_1299_));
 sky130_fd_sc_hs__inv_1 _6333_ (.A(_3786_),
    .Y(_1300_));
 sky130_fd_sc_hs__o21ba_2 _6334_ (.A1(_1300_),
    .A2(_1273_),
    .B1_N(_3785_),
    .X(_1301_));
 sky130_fd_sc_hs__o21bai_2 _6335_ (.A1(_1299_),
    .A2(_1301_),
    .B1_N(_3791_),
    .Y(_1302_));
 sky130_fd_sc_hs__xnor2_4 _6336_ (.A(_1298_),
    .B(_1302_),
    .Y(_1303_));
 sky130_fd_sc_hs__nand2_1 _6337_ (.A(_1088_),
    .B(_1303_),
    .Y(_1304_));
 sky130_fd_sc_hs__a21oi_4 _6338_ (.A1(_1297_),
    .A2(_1304_),
    .B1(_1084_),
    .Y(_1305_));
 sky130_fd_sc_hs__a211oi_4 _6339_ (.A1(net124),
    .A2(_1153_),
    .B1(_1154_),
    .C1(_1305_),
    .Y(_1306_));
 sky130_fd_sc_hs__o21ai_4 _6340_ (.A1(_0810_),
    .A2(_1296_),
    .B1(_1306_),
    .Y(_1307_));
 sky130_fd_sc_hs__nor2_1 _6341_ (.A(_0433_),
    .B(_1290_),
    .Y(_1308_));
 sky130_fd_sc_hs__o21a_1 _6342_ (.A1(_0582_),
    .A2(_1115_),
    .B1(_1116_),
    .X(_1309_));
 sky130_fd_sc_hs__o32a_1 _6343_ (.A1(_1295_),
    .A2(_1307_),
    .A3(_1308_),
    .B1(_1309_),
    .B2(_1305_),
    .X(net295));
 sky130_fd_sc_hs__mux2i_4 _6344_ (.A0(_0584_),
    .A1(net195),
    .S(_1127_),
    .Y(_1310_));
 sky130_fd_sc_hs__nor2_1 _6345_ (.A(_1210_),
    .B(_1310_),
    .Y(_1311_));
 sky130_fd_sc_hs__a31oi_4 _6346_ (.A1(_0095_),
    .A2(_1126_),
    .A3(_0945_),
    .B1(_1311_),
    .Y(_1312_));
 sky130_fd_sc_hs__or2_1 _6347_ (.A(_3792_),
    .B(_3791_),
    .X(_1313_));
 sky130_fd_sc_hs__a21oi_2 _6348_ (.A1(_3801_),
    .A2(_1313_),
    .B1(_3800_),
    .Y(_1314_));
 sky130_fd_sc_hs__inv_1 _6349_ (.A(_1314_),
    .Y(_1315_));
 sky130_fd_sc_hs__a2111o_4 _6350_ (.A1(_3786_),
    .A2(_1280_),
    .B1(_3800_),
    .C1(_3791_),
    .D1(_3785_),
    .X(_1316_));
 sky130_fd_sc_hs__nand2_2 _6351_ (.A(_1315_),
    .B(_1316_),
    .Y(_1317_));
 sky130_fd_sc_hs__xor2_4 _6352_ (.A(_3806_),
    .B(_1317_),
    .X(_1318_));
 sky130_fd_sc_hs__nand2_1 _6353_ (.A(_1147_),
    .B(_1318_),
    .Y(_1319_));
 sky130_fd_sc_hs__clkbuf_16 _6354_ (.A(_1119_),
    .X(_1320_));
 sky130_fd_sc_hs__o211ai_4 _6355_ (.A1(_0584_),
    .A2(_1147_),
    .B1(_1319_),
    .C1(_1320_),
    .Y(_1321_));
 sky130_fd_sc_hs__nor2_2 _6356_ (.A(net125),
    .B(_1125_),
    .Y(_1322_));
 sky130_fd_sc_hs__a21oi_4 _6357_ (.A1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[13] ),
    .A2(_1229_),
    .B1(_1153_),
    .Y(_1323_));
 sky130_fd_sc_hs__nor2_1 _6358_ (.A(_0374_),
    .B(_1191_),
    .Y(_1324_));
 sky130_fd_sc_hs__a21oi_2 _6359_ (.A1(_0584_),
    .A2(_1192_),
    .B1(_1324_),
    .Y(_1325_));
 sky130_fd_sc_hs__o221ai_4 _6360_ (.A1(_1322_),
    .A2(_1323_),
    .B1(_1325_),
    .B2(_1109_),
    .C1(_1231_),
    .Y(_1326_));
 sky130_fd_sc_hs__nor2_1 _6361_ (.A(_0433_),
    .B(_1293_),
    .Y(_1327_));
 sky130_fd_sc_hs__buf_8 _6362_ (.A(_1241_),
    .X(_1328_));
 sky130_fd_sc_hs__o221ai_2 _6363_ (.A1(_0584_),
    .A2(_1122_),
    .B1(_1326_),
    .B2(_1327_),
    .C1(_1328_),
    .Y(_1329_));
 sky130_fd_sc_hs__o211ai_4 _6364_ (.A1(_1082_),
    .A2(_1312_),
    .B1(_1321_),
    .C1(_1329_),
    .Y(net296));
 sky130_fd_sc_hs__a21oi_2 _6365_ (.A1(_0938_),
    .A2(_0945_),
    .B1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[14] ),
    .Y(_1330_));
 sky130_fd_sc_hs__mux2_1 _6366_ (.A0(_0585_),
    .A1(net196),
    .S(_0958_),
    .X(_1331_));
 sky130_fd_sc_hs__o21ai_1 _6367_ (.A1(_1125_),
    .A2(_1331_),
    .B1(_1247_),
    .Y(_1332_));
 sky130_fd_sc_hs__a21oi_1 _6368_ (.A1(_1126_),
    .A2(_1330_),
    .B1(_1332_),
    .Y(_1333_));
 sky130_fd_sc_hs__nand2_1 _6369_ (.A(_0585_),
    .B(_1144_),
    .Y(_1334_));
 sky130_fd_sc_hs__a21oi_2 _6370_ (.A1(_3801_),
    .A2(_3791_),
    .B1(_3800_),
    .Y(_1335_));
 sky130_fd_sc_hs__o31ai_2 _6371_ (.A1(_1299_),
    .A2(_1298_),
    .A3(_1301_),
    .B1(_1335_),
    .Y(_1336_));
 sky130_fd_sc_hs__a21oi_4 _6372_ (.A1(_3806_),
    .A2(_1336_),
    .B1(_3805_),
    .Y(_1337_));
 sky130_fd_sc_hs__xnor2_4 _6373_ (.A(_3813_),
    .B(_1337_),
    .Y(_1338_));
 sky130_fd_sc_hs__nand2_1 _6374_ (.A(_1089_),
    .B(_1338_),
    .Y(_1339_));
 sky130_fd_sc_hs__a21oi_4 _6375_ (.A1(_1334_),
    .A2(_1339_),
    .B1(_1086_),
    .Y(_1340_));
 sky130_fd_sc_hs__nand2b_1 _6376_ (.A_N(_1310_),
    .B(_1264_),
    .Y(_1341_));
 sky130_fd_sc_hs__mux2_1 _6377_ (.A0(_0585_),
    .A1(net16),
    .S(_1107_),
    .X(_1342_));
 sky130_fd_sc_hs__a221oi_4 _6378_ (.A1(net126),
    .A2(_1164_),
    .B1(_1342_),
    .B2(_0430_),
    .C1(_1132_),
    .Y(_1343_));
 sky130_fd_sc_hs__o21ai_1 _6379_ (.A1(_0585_),
    .A2(_1115_),
    .B1(_1116_),
    .Y(_1344_));
 sky130_fd_sc_hs__a21oi_1 _6380_ (.A1(_1341_),
    .A2(_1343_),
    .B1(_1344_),
    .Y(_1345_));
 sky130_fd_sc_hs__or3_1 _6381_ (.A(_1333_),
    .B(_1340_),
    .C(_1345_),
    .X(net297));
 sky130_fd_sc_hs__o21ai_1 _6382_ (.A1(net107),
    .A2(_1122_),
    .B1(_1123_),
    .Y(_1346_));
 sky130_fd_sc_hs__a211oi_2 _6383_ (.A1(_0941_),
    .A2(_0945_),
    .B1(_1079_),
    .C1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[15] ),
    .Y(_1347_));
 sky130_fd_sc_hs__mux2_1 _6384_ (.A0(net107),
    .A1(net197),
    .S(_1211_),
    .X(_1348_));
 sky130_fd_sc_hs__o21ai_1 _6385_ (.A1(_1210_),
    .A2(_1348_),
    .B1(_0386_),
    .Y(_1349_));
 sky130_fd_sc_hs__inv_2 _6386_ (.A(net107),
    .Y(_1350_));
 sky130_fd_sc_hs__nor2_1 _6387_ (.A(_1350_),
    .B(_1107_),
    .Y(_1351_));
 sky130_fd_sc_hs__a21oi_2 _6388_ (.A1(net15),
    .A2(_1151_),
    .B1(_1351_),
    .Y(_1352_));
 sky130_fd_sc_hs__a21oi_2 _6389_ (.A1(net127),
    .A2(_1153_),
    .B1(_1111_),
    .Y(_1353_));
 sky130_fd_sc_hs__o21ai_4 _6390_ (.A1(_1109_),
    .A2(_1352_),
    .B1(_1353_),
    .Y(_1354_));
 sky130_fd_sc_hs__a21oi_1 _6391_ (.A1(_1264_),
    .A2(_1331_),
    .B1(_1354_),
    .Y(_1355_));
 sky130_fd_sc_hs__o21a_1 _6392_ (.A1(_1347_),
    .A2(_1349_),
    .B1(_1355_),
    .X(_1356_));
 sky130_fd_sc_hs__a31o_1 _6393_ (.A1(_3806_),
    .A2(_1315_),
    .A3(_1316_),
    .B1(_3805_),
    .X(_1357_));
 sky130_fd_sc_hs__a21oi_4 _6394_ (.A1(_3813_),
    .A2(_1357_),
    .B1(_3812_),
    .Y(_1358_));
 sky130_fd_sc_hs__xnor2_4 _6395_ (.A(_3824_),
    .B(_1358_),
    .Y(_1359_));
 sky130_fd_sc_hs__nand2_1 _6396_ (.A(_1147_),
    .B(_1359_),
    .Y(_1360_));
 sky130_fd_sc_hs__o21ai_2 _6397_ (.A1(_1350_),
    .A2(_1147_),
    .B1(_1360_),
    .Y(_1361_));
 sky130_fd_sc_hs__nand2_8 _6398_ (.A(_1320_),
    .B(_1361_),
    .Y(_1362_));
 sky130_fd_sc_hs__o21ai_4 _6399_ (.A1(_1346_),
    .A2(_1356_),
    .B1(_1362_),
    .Y(net298));
 sky130_fd_sc_hs__nand2_1 _6400_ (.A(_0814_),
    .B(net108),
    .Y(_1363_));
 sky130_fd_sc_hs__nand2b_1 _6401_ (.A_N(net179),
    .B(_0992_),
    .Y(_1364_));
 sky130_fd_sc_hs__o211ai_2 _6402_ (.A1(net217),
    .A2(_0993_),
    .B1(_1364_),
    .C1(_1037_),
    .Y(_1365_));
 sky130_fd_sc_hs__a21oi_4 _6403_ (.A1(_1363_),
    .A2(_1365_),
    .B1(_0109_),
    .Y(net299));
 sky130_fd_sc_hs__mux2i_4 _6404_ (.A0(_0436_),
    .A1(net198),
    .S(_1127_),
    .Y(_1366_));
 sky130_fd_sc_hs__a311oi_4 _6405_ (.A1(_0920_),
    .A2(_0933_),
    .A3(_0951_),
    .B1(_1076_),
    .C1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[16] ),
    .Y(_1367_));
 sky130_fd_sc_hs__a211oi_1 _6406_ (.A1(_1129_),
    .A2(_1366_),
    .B1(_1367_),
    .C1(_1081_),
    .Y(_1368_));
 sky130_fd_sc_hs__nand2_1 _6407_ (.A(_1264_),
    .B(_1348_),
    .Y(_1369_));
 sky130_fd_sc_hs__mux2_1 _6408_ (.A0(_0436_),
    .A1(net198),
    .S(_1107_),
    .X(_1370_));
 sky130_fd_sc_hs__a221oi_4 _6409_ (.A1(net128),
    .A2(_1164_),
    .B1(_1370_),
    .B2(_0430_),
    .C1(_1132_),
    .Y(_1371_));
 sky130_fd_sc_hs__o21ai_1 _6410_ (.A1(_0436_),
    .A2(_1231_),
    .B1(_1241_),
    .Y(_1372_));
 sky130_fd_sc_hs__a21oi_1 _6411_ (.A1(_1369_),
    .A2(_1371_),
    .B1(_1372_),
    .Y(_1373_));
 sky130_fd_sc_hs__inv_1 _6412_ (.A(_3813_),
    .Y(_1374_));
 sky130_fd_sc_hs__o21bai_1 _6413_ (.A1(_1374_),
    .A2(_1337_),
    .B1_N(_3812_),
    .Y(_1375_));
 sky130_fd_sc_hs__a21oi_4 _6414_ (.A1(_3824_),
    .A2(_1375_),
    .B1(_3823_),
    .Y(_1376_));
 sky130_fd_sc_hs__xor2_4 _6415_ (.A(_3828_),
    .B(_1376_),
    .X(_1377_));
 sky130_fd_sc_hs__nand2_8 _6416_ (.A(_1119_),
    .B(_1146_),
    .Y(_1378_));
 sky130_fd_sc_hs__nand2_1 _6417_ (.A(_3701_),
    .B(_1119_),
    .Y(_1379_));
 sky130_fd_sc_hs__o22ai_4 _6418_ (.A1(_1377_),
    .A2(_1378_),
    .B1(_1379_),
    .B2(_1147_),
    .Y(_1380_));
 sky130_fd_sc_hs__or3_2 _6419_ (.A(_1368_),
    .B(_1373_),
    .C(_1380_),
    .X(net300));
 sky130_fd_sc_hs__a211oi_4 _6420_ (.A1(_0095_),
    .A2(_0954_),
    .B1(_1077_),
    .C1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[17] ),
    .Y(_1381_));
 sky130_fd_sc_hs__mux2_1 _6421_ (.A0(_0446_),
    .A1(net199),
    .S(_1127_),
    .X(_1382_));
 sky130_fd_sc_hs__o21ai_1 _6422_ (.A1(_1126_),
    .A2(_1382_),
    .B1(_1247_),
    .Y(_1383_));
 sky130_fd_sc_hs__inv_1 _6423_ (.A(_3834_),
    .Y(_1384_));
 sky130_fd_sc_hs__nand4_2 _6424_ (.A(_3806_),
    .B(_3813_),
    .C(_3824_),
    .D(_3828_),
    .Y(_1385_));
 sky130_fd_sc_hs__nor2_4 _6425_ (.A(_1314_),
    .B(_1385_),
    .Y(_1386_));
 sky130_fd_sc_hs__inv_1 _6426_ (.A(_3824_),
    .Y(_1387_));
 sky130_fd_sc_hs__a21oi_1 _6427_ (.A1(_3813_),
    .A2(_3805_),
    .B1(_3812_),
    .Y(_1388_));
 sky130_fd_sc_hs__o21bai_2 _6428_ (.A1(_1387_),
    .A2(_1388_),
    .B1_N(_3823_),
    .Y(_1389_));
 sky130_fd_sc_hs__a21oi_2 _6429_ (.A1(_3828_),
    .A2(_1389_),
    .B1(_3827_),
    .Y(_1390_));
 sky130_fd_sc_hs__inv_1 _6430_ (.A(_1390_),
    .Y(_1391_));
 sky130_fd_sc_hs__a21oi_2 _6431_ (.A1(_1316_),
    .A2(_1386_),
    .B1(_1391_),
    .Y(_1392_));
 sky130_fd_sc_hs__xnor2_1 _6432_ (.A(_1384_),
    .B(_1392_),
    .Y(_1393_));
 sky130_fd_sc_hs__nand2_1 _6433_ (.A(_3716_),
    .B(_1178_),
    .Y(_1394_));
 sky130_fd_sc_hs__o21ai_2 _6434_ (.A1(_1178_),
    .A2(_1393_),
    .B1(_1394_),
    .Y(_1395_));
 sky130_fd_sc_hs__nand2_8 _6435_ (.A(_1320_),
    .B(_1395_),
    .Y(_1396_));
 sky130_fd_sc_hs__nor2_1 _6436_ (.A(_0433_),
    .B(_1366_),
    .Y(_1397_));
 sky130_fd_sc_hs__mux2i_2 _6437_ (.A0(_0446_),
    .A1(net199),
    .S(_1134_),
    .Y(_1398_));
 sky130_fd_sc_hs__a21oi_2 _6438_ (.A1(net129),
    .A2(_0123_),
    .B1(_1132_),
    .Y(_1399_));
 sky130_fd_sc_hs__o21ai_2 _6439_ (.A1(_0810_),
    .A2(_1398_),
    .B1(_1399_),
    .Y(_1400_));
 sky130_fd_sc_hs__o221ai_2 _6440_ (.A1(_0446_),
    .A2(_1122_),
    .B1(_1397_),
    .B2(_1400_),
    .C1(_1328_),
    .Y(_1401_));
 sky130_fd_sc_hs__o211ai_4 _6441_ (.A1(_1381_),
    .A2(_1383_),
    .B1(_1396_),
    .C1(_1401_),
    .Y(net301));
 sky130_fd_sc_hs__mux2i_2 _6442_ (.A0(_0449_),
    .A1(net200),
    .S(_1151_),
    .Y(_1402_));
 sky130_fd_sc_hs__a21oi_4 _6443_ (.A1(net130),
    .A2(_0123_),
    .B1(_1132_),
    .Y(_1403_));
 sky130_fd_sc_hs__o21ai_2 _6444_ (.A1(_0810_),
    .A2(_1402_),
    .B1(_1403_),
    .Y(_1404_));
 sky130_fd_sc_hs__a21oi_2 _6445_ (.A1(_0103_),
    .A2(_1382_),
    .B1(_1404_),
    .Y(_1405_));
 sky130_fd_sc_hs__o21ai_1 _6446_ (.A1(_0449_),
    .A2(_1122_),
    .B1(_1123_),
    .Y(_1406_));
 sky130_fd_sc_hs__mux2i_4 _6447_ (.A0(_0449_),
    .A1(net200),
    .S(_1211_),
    .Y(_1407_));
 sky130_fd_sc_hs__nand2_1 _6448_ (.A(_1077_),
    .B(_1407_),
    .Y(_1408_));
 sky130_fd_sc_hs__a311o_1 _6449_ (.A1(_0938_),
    .A2(_0933_),
    .A3(_0951_),
    .B1(_1129_),
    .C1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[18] ),
    .X(_1409_));
 sky130_fd_sc_hs__nand3_1 _6450_ (.A(_1247_),
    .B(_1408_),
    .C(_1409_),
    .Y(_1410_));
 sky130_fd_sc_hs__or2_1 _6451_ (.A(_1298_),
    .B(_1385_),
    .X(_1411_));
 sky130_fd_sc_hs__nor2_1 _6452_ (.A(_1335_),
    .B(_1385_),
    .Y(_1412_));
 sky130_fd_sc_hs__a211oi_4 _6453_ (.A1(_3828_),
    .A2(_1389_),
    .B1(_1412_),
    .C1(_3827_),
    .Y(_1413_));
 sky130_fd_sc_hs__o31ai_4 _6454_ (.A1(_1299_),
    .A2(_1301_),
    .A3(_1411_),
    .B1(_1413_),
    .Y(_1414_));
 sky130_fd_sc_hs__a21oi_1 _6455_ (.A1(_3834_),
    .A2(_1414_),
    .B1(_3833_),
    .Y(_1415_));
 sky130_fd_sc_hs__xnor2_1 _6456_ (.A(_3840_),
    .B(_1415_),
    .Y(_1416_));
 sky130_fd_sc_hs__mux2_2 _6457_ (.A0(_3718_),
    .A1(_1416_),
    .S(_1089_),
    .X(_1417_));
 sky130_fd_sc_hs__nand2_8 _6458_ (.A(_1320_),
    .B(_1417_),
    .Y(_1418_));
 sky130_fd_sc_hs__o211ai_4 _6459_ (.A1(_1405_),
    .A2(_1406_),
    .B1(_1410_),
    .C1(_1418_),
    .Y(net302));
 sky130_fd_sc_hs__or2_1 _6460_ (.A(_0586_),
    .B(_1115_),
    .X(_1419_));
 sky130_fd_sc_hs__inv_2 _6461_ (.A(_3846_),
    .Y(_1420_));
 sky130_fd_sc_hs__o21bai_1 _6462_ (.A1(_1384_),
    .A2(_1392_),
    .B1_N(_3833_),
    .Y(_1421_));
 sky130_fd_sc_hs__a21oi_4 _6463_ (.A1(_3840_),
    .A2(_1421_),
    .B1(_3839_),
    .Y(_1422_));
 sky130_fd_sc_hs__xnor2_4 _6464_ (.A(_1420_),
    .B(_1422_),
    .Y(_1423_));
 sky130_fd_sc_hs__nand2_1 _6465_ (.A(_3726_),
    .B(_1119_),
    .Y(_1424_));
 sky130_fd_sc_hs__o22ai_4 _6466_ (.A1(_1378_),
    .A2(_1423_),
    .B1(_1424_),
    .B2(_1147_),
    .Y(_1425_));
 sky130_fd_sc_hs__a21oi_1 _6467_ (.A1(_1328_),
    .A2(_1419_),
    .B1(_1425_),
    .Y(_1426_));
 sky130_fd_sc_hs__a311o_2 _6468_ (.A1(_0941_),
    .A2(_0933_),
    .A3(_0951_),
    .B1(_1076_),
    .C1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[19] ),
    .X(_1427_));
 sky130_fd_sc_hs__mux2i_4 _6469_ (.A0(_0586_),
    .A1(net201),
    .S(_1211_),
    .Y(_1428_));
 sky130_fd_sc_hs__nand2_1 _6470_ (.A(_1077_),
    .B(_1428_),
    .Y(_1429_));
 sky130_fd_sc_hs__mux2i_4 _6471_ (.A0(_0586_),
    .A1(net201),
    .S(_1151_),
    .Y(_1430_));
 sky130_fd_sc_hs__a21oi_4 _6472_ (.A1(net131),
    .A2(_1164_),
    .B1(_1154_),
    .Y(_1431_));
 sky130_fd_sc_hs__o221ai_4 _6473_ (.A1(_0391_),
    .A2(_1407_),
    .B1(_1430_),
    .B2(_1109_),
    .C1(_1431_),
    .Y(_1432_));
 sky130_fd_sc_hs__a311oi_4 _6474_ (.A1(_0386_),
    .A2(_1427_),
    .A3(_1429_),
    .B1(_1432_),
    .C1(_1425_),
    .Y(_1433_));
 sky130_fd_sc_hs__nor2_4 _6475_ (.A(_1426_),
    .B(_1433_),
    .Y(net303));
 sky130_fd_sc_hs__a311oi_2 _6476_ (.A1(_0920_),
    .A2(_0933_),
    .A3(_0962_),
    .B1(_1079_),
    .C1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[20] ),
    .Y(_1434_));
 sky130_fd_sc_hs__mux2_1 _6477_ (.A0(_0588_),
    .A1(net203),
    .S(_1211_),
    .X(_1435_));
 sky130_fd_sc_hs__nor2_1 _6478_ (.A(_1210_),
    .B(_1435_),
    .Y(_1436_));
 sky130_fd_sc_hs__nor3_1 _6479_ (.A(_1081_),
    .B(_1434_),
    .C(_1436_),
    .Y(_1437_));
 sky130_fd_sc_hs__nand2b_1 _6480_ (.A_N(_1428_),
    .B(_0102_),
    .Y(_1438_));
 sky130_fd_sc_hs__mux2_1 _6481_ (.A0(_0588_),
    .A1(net203),
    .S(_1107_),
    .X(_1439_));
 sky130_fd_sc_hs__a221oi_4 _6482_ (.A1(net133),
    .A2(_1164_),
    .B1(_1439_),
    .B2(_0430_),
    .C1(_1154_),
    .Y(_1440_));
 sky130_fd_sc_hs__o21ai_1 _6483_ (.A1(_0588_),
    .A2(_1114_),
    .B1(_1241_),
    .Y(_1441_));
 sky130_fd_sc_hs__a21oi_1 _6484_ (.A1(_1438_),
    .A2(_1440_),
    .B1(_1441_),
    .Y(_1442_));
 sky130_fd_sc_hs__nand2_1 _6485_ (.A(_3730_),
    .B(_1144_),
    .Y(_1443_));
 sky130_fd_sc_hs__nand2_1 _6486_ (.A(_3840_),
    .B(_3833_),
    .Y(_1444_));
 sky130_fd_sc_hs__clkinv_1 _6487_ (.A(_1444_),
    .Y(_1445_));
 sky130_fd_sc_hs__a311oi_4 _6488_ (.A1(_3834_),
    .A2(_3840_),
    .A3(_1414_),
    .B1(_1445_),
    .C1(_3839_),
    .Y(_1446_));
 sky130_fd_sc_hs__o21bai_2 _6489_ (.A1(_1420_),
    .A2(_1446_),
    .B1_N(_3845_),
    .Y(_1447_));
 sky130_fd_sc_hs__xor2_4 _6490_ (.A(_3852_),
    .B(_1447_),
    .X(_1448_));
 sky130_fd_sc_hs__nand2_1 _6491_ (.A(_1147_),
    .B(_1448_),
    .Y(_1449_));
 sky130_fd_sc_hs__a21oi_4 _6492_ (.A1(_1443_),
    .A2(_1449_),
    .B1(_1086_),
    .Y(_1450_));
 sky130_fd_sc_hs__or3_1 _6493_ (.A(_1437_),
    .B(_1442_),
    .C(_1450_),
    .X(net304));
 sky130_fd_sc_hs__mux2_1 _6494_ (.A0(net109),
    .A1(net204),
    .S(_1211_),
    .X(_1451_));
 sky130_fd_sc_hs__nor2_2 _6495_ (.A(_1126_),
    .B(_1451_),
    .Y(_1452_));
 sky130_fd_sc_hs__a211oi_4 _6496_ (.A1(_0095_),
    .A2(_0964_),
    .B1(_1077_),
    .C1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[21] ),
    .Y(_1453_));
 sky130_fd_sc_hs__nand3_1 _6497_ (.A(_3858_),
    .B(_1119_),
    .C(_1146_),
    .Y(_1454_));
 sky130_fd_sc_hs__nand3b_4 _6498_ (.A_N(_3858_),
    .B(_1119_),
    .C(_1089_),
    .Y(_1455_));
 sky130_fd_sc_hs__nand2_1 _6499_ (.A(_3846_),
    .B(_3852_),
    .Y(_1456_));
 sky130_fd_sc_hs__a21o_1 _6500_ (.A1(_3852_),
    .A2(_3845_),
    .B1(_3851_),
    .X(_1457_));
 sky130_fd_sc_hs__o21bai_4 _6501_ (.A1(_1422_),
    .A2(_1456_),
    .B1_N(_1457_),
    .Y(_1458_));
 sky130_fd_sc_hs__mux2i_4 _6502_ (.A0(_1454_),
    .A1(_1455_),
    .S(_1458_),
    .Y(_1459_));
 sky130_fd_sc_hs__a31oi_4 _6503_ (.A1(_3739_),
    .A2(_1320_),
    .A3(_1178_),
    .B1(_1459_),
    .Y(_1460_));
 sky130_fd_sc_hs__and2_1 _6504_ (.A(_0103_),
    .B(_1435_),
    .X(_1461_));
 sky130_fd_sc_hs__a21oi_4 _6505_ (.A1(net134),
    .A2(_0122_),
    .B1(_1111_),
    .Y(_1462_));
 sky130_fd_sc_hs__o21ai_1 _6506_ (.A1(net204),
    .A2(_1192_),
    .B1(_0430_),
    .Y(_1463_));
 sky130_fd_sc_hs__nand2_1 _6507_ (.A(_1192_),
    .B(_1462_),
    .Y(_1464_));
 sky130_fd_sc_hs__a21oi_2 _6508_ (.A1(_1114_),
    .A2(_1464_),
    .B1(net109),
    .Y(_1465_));
 sky130_fd_sc_hs__a21oi_4 _6509_ (.A1(_1462_),
    .A2(_1463_),
    .B1(_1465_),
    .Y(_1466_));
 sky130_fd_sc_hs__o21ai_1 _6510_ (.A1(_1461_),
    .A2(_1466_),
    .B1(_1242_),
    .Y(_1467_));
 sky130_fd_sc_hs__o311ai_4 _6511_ (.A1(_1082_),
    .A2(_1452_),
    .A3(_1453_),
    .B1(_1460_),
    .C1(_1467_),
    .Y(net305));
 sky130_fd_sc_hs__mux2i_4 _6512_ (.A0(_0520_),
    .A1(net205),
    .S(_1127_),
    .Y(_1468_));
 sky130_fd_sc_hs__nand2_1 _6513_ (.A(_1077_),
    .B(_1468_),
    .Y(_1469_));
 sky130_fd_sc_hs__a311o_1 _6514_ (.A1(_0938_),
    .A2(_0933_),
    .A3(_0962_),
    .B1(_1079_),
    .C1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[22] ),
    .X(_1470_));
 sky130_fd_sc_hs__nand3_2 _6515_ (.A(_3846_),
    .B(_3852_),
    .C(_3858_),
    .Y(_1471_));
 sky130_fd_sc_hs__a21oi_4 _6516_ (.A1(_3858_),
    .A2(_1457_),
    .B1(_3857_),
    .Y(_1472_));
 sky130_fd_sc_hs__o21ai_1 _6517_ (.A1(_1446_),
    .A2(_1471_),
    .B1(_1472_),
    .Y(_1473_));
 sky130_fd_sc_hs__xnor2_2 _6518_ (.A(_3864_),
    .B(_1473_),
    .Y(_1474_));
 sky130_fd_sc_hs__nand2_1 _6519_ (.A(_3749_),
    .B(_1143_),
    .Y(_1475_));
 sky130_fd_sc_hs__o21ai_1 _6520_ (.A1(_1143_),
    .A2(_1474_),
    .B1(_1475_),
    .Y(_1476_));
 sky130_fd_sc_hs__and2_4 _6521_ (.A(_1320_),
    .B(_1476_),
    .X(_1477_));
 sky130_fd_sc_hs__nand2_1 _6522_ (.A(_1264_),
    .B(_1451_),
    .Y(_1478_));
 sky130_fd_sc_hs__mux2_1 _6523_ (.A0(_0520_),
    .A1(net205),
    .S(_1106_),
    .X(_1479_));
 sky130_fd_sc_hs__a221oi_4 _6524_ (.A1(net135),
    .A2(_1164_),
    .B1(_1479_),
    .B2(_0378_),
    .C1(_1154_),
    .Y(_1480_));
 sky130_fd_sc_hs__o21ai_1 _6525_ (.A1(_0520_),
    .A2(_1114_),
    .B1(_1241_),
    .Y(_1481_));
 sky130_fd_sc_hs__a21oi_1 _6526_ (.A1(_1478_),
    .A2(_1480_),
    .B1(_1481_),
    .Y(_1482_));
 sky130_fd_sc_hs__a311o_1 _6527_ (.A1(_1247_),
    .A2(_1469_),
    .A3(_1470_),
    .B1(_1477_),
    .C1(_1482_),
    .X(net306));
 sky130_fd_sc_hs__mux2_1 _6528_ (.A0(_0526_),
    .A1(net206),
    .S(_1211_),
    .X(_1483_));
 sky130_fd_sc_hs__nand2_1 _6529_ (.A(_1129_),
    .B(_1483_),
    .Y(_1484_));
 sky130_fd_sc_hs__nand4_1 _6530_ (.A(_0941_),
    .B(_1125_),
    .C(_0933_),
    .D(_0962_),
    .Y(_1485_));
 sky130_fd_sc_hs__a21oi_1 _6531_ (.A1(_1484_),
    .A2(_1485_),
    .B1(_1082_),
    .Y(_1486_));
 sky130_fd_sc_hs__nand2_1 _6532_ (.A(_2347_),
    .B(_1144_),
    .Y(_1487_));
 sky130_fd_sc_hs__inv_1 _6533_ (.A(_3864_),
    .Y(_1488_));
 sky130_fd_sc_hs__or2_1 _6534_ (.A(_3834_),
    .B(_3833_),
    .X(_1489_));
 sky130_fd_sc_hs__a21oi_1 _6535_ (.A1(_3840_),
    .A2(_1489_),
    .B1(_3839_),
    .Y(_1490_));
 sky130_fd_sc_hs__o21a_1 _6536_ (.A1(_1471_),
    .A2(_1490_),
    .B1(_1472_),
    .X(_1491_));
 sky130_fd_sc_hs__nor2_1 _6537_ (.A(_3833_),
    .B(_3839_),
    .Y(_1492_));
 sky130_fd_sc_hs__nand3_1 _6538_ (.A(_1390_),
    .B(_1472_),
    .C(_1492_),
    .Y(_1493_));
 sky130_fd_sc_hs__a21oi_4 _6539_ (.A1(_1316_),
    .A2(_1386_),
    .B1(_1493_),
    .Y(_1494_));
 sky130_fd_sc_hs__nor3_1 _6540_ (.A(_1488_),
    .B(_1491_),
    .C(_1494_),
    .Y(_1495_));
 sky130_fd_sc_hs__nor2_1 _6541_ (.A(_3863_),
    .B(_1495_),
    .Y(_1496_));
 sky130_fd_sc_hs__xnor2_1 _6542_ (.A(_3870_),
    .B(_1496_),
    .Y(_1497_));
 sky130_fd_sc_hs__nand2_2 _6543_ (.A(_1089_),
    .B(_1497_),
    .Y(_1498_));
 sky130_fd_sc_hs__a21oi_4 _6544_ (.A1(_1487_),
    .A2(_1498_),
    .B1(_1086_),
    .Y(_1499_));
 sky130_fd_sc_hs__nor2_4 _6545_ (.A(net136),
    .B(_0818_),
    .Y(_1500_));
 sky130_fd_sc_hs__a21oi_1 _6546_ (.A1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[23] ),
    .A2(_1229_),
    .B1(_0122_),
    .Y(_1501_));
 sky130_fd_sc_hs__mux2i_1 _6547_ (.A0(_0526_),
    .A1(net206),
    .S(_1107_),
    .Y(_1502_));
 sky130_fd_sc_hs__o221a_1 _6548_ (.A1(_1500_),
    .A2(_1501_),
    .B1(_1502_),
    .B2(_1109_),
    .C1(_1114_),
    .X(_1503_));
 sky130_fd_sc_hs__nand2b_1 _6549_ (.A_N(_1468_),
    .B(_1264_),
    .Y(_1504_));
 sky130_fd_sc_hs__o21ai_1 _6550_ (.A1(_0526_),
    .A2(_1231_),
    .B1(_1116_),
    .Y(_1505_));
 sky130_fd_sc_hs__a21oi_1 _6551_ (.A1(_1503_),
    .A2(_1504_),
    .B1(_1505_),
    .Y(_1506_));
 sky130_fd_sc_hs__or3_2 _6552_ (.A(_1486_),
    .B(_1499_),
    .C(_1506_),
    .X(net307));
 sky130_fd_sc_hs__mux2i_4 _6553_ (.A0(_0527_),
    .A1(net13),
    .S(_1211_),
    .Y(_1507_));
 sky130_fd_sc_hs__a211oi_1 _6554_ (.A1(_0920_),
    .A2(_0969_),
    .B1(_1076_),
    .C1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[24] ),
    .Y(_1508_));
 sky130_fd_sc_hs__a211oi_1 _6555_ (.A1(_1129_),
    .A2(_1507_),
    .B1(_1508_),
    .C1(_1081_),
    .Y(_1509_));
 sky130_fd_sc_hs__nand2b_1 _6556_ (.A_N(_3839_),
    .B(_1472_),
    .Y(_1510_));
 sky130_fd_sc_hs__a311o_1 _6557_ (.A1(_3834_),
    .A2(_3840_),
    .A3(_1414_),
    .B1(_1445_),
    .C1(_1510_),
    .X(_1511_));
 sky130_fd_sc_hs__a21oi_2 _6558_ (.A1(_1471_),
    .A2(_1472_),
    .B1(_1488_),
    .Y(_1512_));
 sky130_fd_sc_hs__a21oi_1 _6559_ (.A1(_1511_),
    .A2(_1512_),
    .B1(_3863_),
    .Y(_1513_));
 sky130_fd_sc_hs__nor2b_1 _6560_ (.A(_1513_),
    .B_N(_3870_),
    .Y(_1514_));
 sky130_fd_sc_hs__nor2_1 _6561_ (.A(_3869_),
    .B(_1514_),
    .Y(_1515_));
 sky130_fd_sc_hs__or4_1 _6562_ (.A(_3876_),
    .B(_1084_),
    .C(_1143_),
    .D(_1515_),
    .X(_1516_));
 sky130_fd_sc_hs__nand4_1 _6563_ (.A(_3876_),
    .B(_1119_),
    .C(_1146_),
    .D(_1515_),
    .Y(_1517_));
 sky130_fd_sc_hs__o311ai_2 _6564_ (.A1(_1085_),
    .A2(_1146_),
    .A3(_1232_),
    .B1(_1516_),
    .C1(_1517_),
    .Y(_1518_));
 sky130_fd_sc_hs__nand2_1 _6565_ (.A(_0527_),
    .B(_1192_),
    .Y(_1519_));
 sky130_fd_sc_hs__nand2_1 _6566_ (.A(net13),
    .B(_1134_),
    .Y(_1520_));
 sky130_fd_sc_hs__nand2_1 _6567_ (.A(_0105_),
    .B(_0430_),
    .Y(_1521_));
 sky130_fd_sc_hs__a21oi_1 _6568_ (.A1(_1519_),
    .A2(_1520_),
    .B1(_1521_),
    .Y(_1522_));
 sky130_fd_sc_hs__nand2_1 _6569_ (.A(_1264_),
    .B(_1483_),
    .Y(_1523_));
 sky130_fd_sc_hs__a21oi_4 _6570_ (.A1(net137),
    .A2(_0123_),
    .B1(_1132_),
    .Y(_1524_));
 sky130_fd_sc_hs__o21ai_1 _6571_ (.A1(_0527_),
    .A2(_1231_),
    .B1(_1241_),
    .Y(_1525_));
 sky130_fd_sc_hs__a21oi_1 _6572_ (.A1(_1523_),
    .A2(_1524_),
    .B1(_1525_),
    .Y(_1526_));
 sky130_fd_sc_hs__or4_1 _6573_ (.A(_1509_),
    .B(_1518_),
    .C(_1522_),
    .D(_1526_),
    .X(net308));
 sky130_fd_sc_hs__a21oi_1 _6574_ (.A1(_0095_),
    .A2(_0969_),
    .B1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[25] ),
    .Y(_1527_));
 sky130_fd_sc_hs__mux2_1 _6575_ (.A0(_0529_),
    .A1(net208),
    .S(_0958_),
    .X(_1528_));
 sky130_fd_sc_hs__o21ai_1 _6576_ (.A1(_1125_),
    .A2(_1528_),
    .B1(_1247_),
    .Y(_1529_));
 sky130_fd_sc_hs__a21oi_1 _6577_ (.A1(_1210_),
    .A2(_1527_),
    .B1(_1529_),
    .Y(_1530_));
 sky130_fd_sc_hs__nand2_1 _6578_ (.A(_1144_),
    .B(_1253_),
    .Y(_1531_));
 sky130_fd_sc_hs__o21a_1 _6579_ (.A1(_3864_),
    .A2(_3863_),
    .B1(_3870_),
    .X(_1532_));
 sky130_fd_sc_hs__o21ai_1 _6580_ (.A1(_3869_),
    .A2(_1532_),
    .B1(_3876_),
    .Y(_1533_));
 sky130_fd_sc_hs__nor2_1 _6581_ (.A(_3863_),
    .B(_3869_),
    .Y(_1534_));
 sky130_fd_sc_hs__o21a_1 _6582_ (.A1(_1491_),
    .A2(_1494_),
    .B1(_1534_),
    .X(_1535_));
 sky130_fd_sc_hs__o21bai_1 _6583_ (.A1(_1533_),
    .A2(_1535_),
    .B1_N(_3875_),
    .Y(_1536_));
 sky130_fd_sc_hs__xor2_1 _6584_ (.A(_3882_),
    .B(_1536_),
    .X(_1537_));
 sky130_fd_sc_hs__nand2_2 _6585_ (.A(_1089_),
    .B(_1537_),
    .Y(_1538_));
 sky130_fd_sc_hs__a21oi_4 _6586_ (.A1(_1531_),
    .A2(_1538_),
    .B1(_1086_),
    .Y(_1539_));
 sky130_fd_sc_hs__nor2_1 _6587_ (.A(_0391_),
    .B(_1507_),
    .Y(_1540_));
 sky130_fd_sc_hs__mux2i_1 _6588_ (.A0(_0529_),
    .A1(net208),
    .S(_1107_),
    .Y(_1541_));
 sky130_fd_sc_hs__a21oi_2 _6589_ (.A1(net138),
    .A2(_1153_),
    .B1(_1111_),
    .Y(_1542_));
 sky130_fd_sc_hs__o21ai_1 _6590_ (.A1(_1109_),
    .A2(_1541_),
    .B1(_1542_),
    .Y(_1543_));
 sky130_fd_sc_hs__o221a_1 _6591_ (.A1(_0529_),
    .A2(_1114_),
    .B1(_1540_),
    .B2(_1543_),
    .C1(_1116_),
    .X(_1544_));
 sky130_fd_sc_hs__or3_1 _6592_ (.A(_1530_),
    .B(_1539_),
    .C(_1544_),
    .X(net309));
 sky130_fd_sc_hs__nor2_1 _6593_ (.A(_0317_),
    .B(_1035_),
    .Y(_1545_));
 sky130_fd_sc_hs__a21oi_2 _6594_ (.A1(net180),
    .A2(_1035_),
    .B1(_1545_),
    .Y(_1546_));
 sky130_fd_sc_hs__nor2_1 _6595_ (.A(_0995_),
    .B(net110),
    .Y(_1547_));
 sky130_fd_sc_hs__a211oi_4 _6596_ (.A1(_0091_),
    .A2(_1546_),
    .B1(_1547_),
    .C1(_0788_),
    .Y(net310));
 sky130_fd_sc_hs__mux2_2 _6597_ (.A0(_0565_),
    .A1(net209),
    .S(_0959_),
    .X(_1548_));
 sky130_fd_sc_hs__a211o_1 _6598_ (.A1(_0938_),
    .A2(_0969_),
    .B1(_1129_),
    .C1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[26] ),
    .X(_1549_));
 sky130_fd_sc_hs__o211ai_4 _6599_ (.A1(_1126_),
    .A2(_1548_),
    .B1(_1549_),
    .C1(_1247_),
    .Y(_1550_));
 sky130_fd_sc_hs__nor3_1 _6600_ (.A(_3888_),
    .B(_1084_),
    .C(_1143_),
    .Y(_1551_));
 sky130_fd_sc_hs__nor4b_1 _6601_ (.A(_3881_),
    .B(_1084_),
    .C(_1143_),
    .D_N(_3888_),
    .Y(_1552_));
 sky130_fd_sc_hs__o21a_1 _6602_ (.A1(_3876_),
    .A2(_3875_),
    .B1(_3882_),
    .X(_1553_));
 sky130_fd_sc_hs__o31ai_1 _6603_ (.A1(_3869_),
    .A2(_3875_),
    .A3(_1514_),
    .B1(_1553_),
    .Y(_1554_));
 sky130_fd_sc_hs__mux2_1 _6604_ (.A0(_1551_),
    .A1(_1552_),
    .S(_1554_),
    .X(_1555_));
 sky130_fd_sc_hs__nor4b_2 _6605_ (.A(_3888_),
    .B(_1144_),
    .C(_1085_),
    .D_N(_3881_),
    .Y(_1556_));
 sky130_fd_sc_hs__a311oi_4 _6606_ (.A1(_1320_),
    .A2(_1178_),
    .A3(_1274_),
    .B1(_1555_),
    .C1(_1556_),
    .Y(_1557_));
 sky130_fd_sc_hs__a21oi_4 _6607_ (.A1(net139),
    .A2(_0123_),
    .B1(_1132_),
    .Y(_1558_));
 sky130_fd_sc_hs__nor4_2 _6608_ (.A(_0381_),
    .B(_0128_),
    .C(_0213_),
    .D(_1191_),
    .Y(_1559_));
 sky130_fd_sc_hs__and4_1 _6609_ (.A(_0378_),
    .B(_0128_),
    .C(_0213_),
    .D(_1107_),
    .X(_1560_));
 sky130_fd_sc_hs__and3_1 _6610_ (.A(_0378_),
    .B(_0565_),
    .C(_1191_),
    .X(_1561_));
 sky130_fd_sc_hs__a2111oi_2 _6611_ (.A1(_1264_),
    .A2(_1528_),
    .B1(_1559_),
    .C1(_1560_),
    .D1(_1561_),
    .Y(_1562_));
 sky130_fd_sc_hs__o21ai_1 _6612_ (.A1(_0565_),
    .A2(_1115_),
    .B1(_1116_),
    .Y(_1563_));
 sky130_fd_sc_hs__a21o_1 _6613_ (.A1(_1558_),
    .A2(_1562_),
    .B1(_1563_),
    .X(_1564_));
 sky130_fd_sc_hs__nand3_4 _6614_ (.A(_1550_),
    .B(_1557_),
    .C(_1564_),
    .Y(net311));
 sky130_fd_sc_hs__mux2i_4 _6615_ (.A0(_0566_),
    .A1(net210),
    .S(_0959_),
    .Y(_1565_));
 sky130_fd_sc_hs__nor2_1 _6616_ (.A(_1210_),
    .B(_1565_),
    .Y(_1566_));
 sky130_fd_sc_hs__a31oi_4 _6617_ (.A1(_0941_),
    .A2(_1126_),
    .A3(_0969_),
    .B1(_1566_),
    .Y(_1567_));
 sky130_fd_sc_hs__nor2_2 _6618_ (.A(_3875_),
    .B(_3881_),
    .Y(_1568_));
 sky130_fd_sc_hs__o211ai_2 _6619_ (.A1(_1491_),
    .A2(_1494_),
    .B1(_1534_),
    .C1(_1568_),
    .Y(_1569_));
 sky130_fd_sc_hs__nor2_1 _6620_ (.A(_3882_),
    .B(_3881_),
    .Y(_1570_));
 sky130_fd_sc_hs__a21oi_2 _6621_ (.A1(_1533_),
    .A2(_1568_),
    .B1(_1570_),
    .Y(_1571_));
 sky130_fd_sc_hs__a31oi_1 _6622_ (.A1(_3888_),
    .A2(_1569_),
    .A3(_1571_),
    .B1(_3887_),
    .Y(_1572_));
 sky130_fd_sc_hs__xnor2_1 _6623_ (.A(_3894_),
    .B(_1572_),
    .Y(_1573_));
 sky130_fd_sc_hs__mux2_2 _6624_ (.A0(_1282_),
    .A1(_1573_),
    .S(_1089_),
    .X(_1574_));
 sky130_fd_sc_hs__nand2_8 _6625_ (.A(_1320_),
    .B(_1574_),
    .Y(_1575_));
 sky130_fd_sc_hs__nand2b_1 _6626_ (.A_N(_0566_),
    .B(_1191_),
    .Y(_1576_));
 sky130_fd_sc_hs__o211ai_1 _6627_ (.A1(net210),
    .A2(_1192_),
    .B1(_1576_),
    .C1(_0430_),
    .Y(_1577_));
 sky130_fd_sc_hs__a21oi_1 _6628_ (.A1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[27] ),
    .A2(_1229_),
    .B1(_1153_),
    .Y(_1578_));
 sky130_fd_sc_hs__o21bai_1 _6629_ (.A1(net140),
    .A2(_1125_),
    .B1_N(_1578_),
    .Y(_1579_));
 sky130_fd_sc_hs__a31oi_2 _6630_ (.A1(_1115_),
    .A2(_1577_),
    .A3(_1579_),
    .B1(_1246_),
    .Y(_1580_));
 sky130_fd_sc_hs__a31oi_2 _6631_ (.A1(_0103_),
    .A2(_1123_),
    .A3(_1548_),
    .B1(_1580_),
    .Y(_1581_));
 sky130_fd_sc_hs__o211ai_4 _6632_ (.A1(_1082_),
    .A2(_1567_),
    .B1(_1575_),
    .C1(_1581_),
    .Y(net312));
 sky130_fd_sc_hs__a311oi_2 _6633_ (.A1(_0920_),
    .A2(_0974_),
    .A3(_0962_),
    .B1(_1129_),
    .C1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[28] ),
    .Y(_1582_));
 sky130_fd_sc_hs__inv_1 _6634_ (.A(net111),
    .Y(_1583_));
 sky130_fd_sc_hs__nor2_1 _6635_ (.A(_1583_),
    .B(_0958_),
    .Y(_1584_));
 sky130_fd_sc_hs__a211oi_1 _6636_ (.A1(net12),
    .A2(_0959_),
    .B1(_1584_),
    .C1(_1210_),
    .Y(_1585_));
 sky130_fd_sc_hs__nor3_1 _6637_ (.A(_1082_),
    .B(_1582_),
    .C(_1585_),
    .Y(_1586_));
 sky130_fd_sc_hs__o21a_1 _6638_ (.A1(_3888_),
    .A2(_3887_),
    .B1(_3894_),
    .X(_1587_));
 sky130_fd_sc_hs__nand4_1 _6639_ (.A(_3870_),
    .B(_3876_),
    .C(_3882_),
    .D(_1587_),
    .Y(_1588_));
 sky130_fd_sc_hs__nand3b_2 _6640_ (.A_N(_1588_),
    .B(_1511_),
    .C(_1512_),
    .Y(_1589_));
 sky130_fd_sc_hs__a21oi_1 _6641_ (.A1(_3876_),
    .A2(_3869_),
    .B1(_3875_),
    .Y(_1590_));
 sky130_fd_sc_hs__nor2b_1 _6642_ (.A(_1590_),
    .B_N(_3882_),
    .Y(_1591_));
 sky130_fd_sc_hs__and4_1 _6643_ (.A(_3870_),
    .B(_3876_),
    .C(_3882_),
    .D(_3863_),
    .X(_1592_));
 sky130_fd_sc_hs__o41ai_1 _6644_ (.A1(_3881_),
    .A2(_3887_),
    .A3(_1591_),
    .A4(_1592_),
    .B1(_1587_),
    .Y(_1593_));
 sky130_fd_sc_hs__nand3b_1 _6645_ (.A_N(_3893_),
    .B(_1589_),
    .C(_1593_),
    .Y(_1594_));
 sky130_fd_sc_hs__xnor2_1 _6646_ (.A(_3900_),
    .B(_1594_),
    .Y(_1595_));
 sky130_fd_sc_hs__nand2_1 _6647_ (.A(_1178_),
    .B(_1303_),
    .Y(_1596_));
 sky130_fd_sc_hs__o21ai_2 _6648_ (.A1(_1178_),
    .A2(_1595_),
    .B1(_1596_),
    .Y(_1597_));
 sky130_fd_sc_hs__nand2_8 _6649_ (.A(_1320_),
    .B(_1597_),
    .Y(_1598_));
 sky130_fd_sc_hs__o21ai_2 _6650_ (.A1(net141),
    .A2(_1125_),
    .B1(_0123_),
    .Y(_1599_));
 sky130_fd_sc_hs__o21ai_1 _6651_ (.A1(_1583_),
    .A2(_1231_),
    .B1(_1599_),
    .Y(_1600_));
 sky130_fd_sc_hs__nor2_1 _6652_ (.A(_0433_),
    .B(_1565_),
    .Y(_1601_));
 sky130_fd_sc_hs__nand2_1 _6653_ (.A(net111),
    .B(_1192_),
    .Y(_1602_));
 sky130_fd_sc_hs__nand2_1 _6654_ (.A(net12),
    .B(_1134_),
    .Y(_1603_));
 sky130_fd_sc_hs__a21oi_1 _6655_ (.A1(_1602_),
    .A2(_1603_),
    .B1(_0810_),
    .Y(_1604_));
 sky130_fd_sc_hs__o31ai_1 _6656_ (.A1(_1600_),
    .A2(_1601_),
    .A3(_1604_),
    .B1(_1242_),
    .Y(_1605_));
 sky130_fd_sc_hs__nand3b_4 _6657_ (.A_N(_1586_),
    .B(_1598_),
    .C(_1605_),
    .Y(net313));
 sky130_fd_sc_hs__buf_8 _6658_ (.A(_1241_),
    .X(_1606_));
 sky130_fd_sc_hs__nand4_1 _6659_ (.A(_0097_),
    .B(_0095_),
    .C(_0958_),
    .D(_0962_),
    .Y(_1607_));
 sky130_fd_sc_hs__nor2_1 _6660_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[29] ),
    .B(_1075_),
    .Y(_1608_));
 sky130_fd_sc_hs__mux2i_4 _6661_ (.A0(net112),
    .A1(net11),
    .S(_0958_),
    .Y(_1609_));
 sky130_fd_sc_hs__a22oi_1 _6662_ (.A1(_1607_),
    .A2(_1608_),
    .B1(_1609_),
    .B2(_1076_),
    .Y(_1610_));
 sky130_fd_sc_hs__inv_1 _6663_ (.A(net112),
    .Y(_1611_));
 sky130_fd_sc_hs__nand2b_1 _6664_ (.A_N(_1110_),
    .B(_1611_),
    .Y(_1612_));
 sky130_fd_sc_hs__nor2_1 _6665_ (.A(_1611_),
    .B(_1106_),
    .Y(_1613_));
 sky130_fd_sc_hs__a21oi_1 _6666_ (.A1(net9),
    .A2(_1107_),
    .B1(_1613_),
    .Y(_1614_));
 sky130_fd_sc_hs__a21oi_2 _6667_ (.A1(net142),
    .A2(_0122_),
    .B1(_1111_),
    .Y(_1615_));
 sky130_fd_sc_hs__o21ai_1 _6668_ (.A1(_0381_),
    .A2(_1614_),
    .B1(_1615_),
    .Y(_1616_));
 sky130_fd_sc_hs__a31o_1 _6669_ (.A1(net12),
    .A2(_1127_),
    .A3(_1612_),
    .B1(_1584_),
    .X(_1617_));
 sky130_fd_sc_hs__a222o_1 _6670_ (.A1(_0386_),
    .A2(_1610_),
    .B1(_1612_),
    .B2(_1616_),
    .C1(_1617_),
    .C2(_1264_),
    .X(_1618_));
 sky130_fd_sc_hs__and3_1 _6671_ (.A(_3888_),
    .B(_3894_),
    .C(_3900_),
    .X(_1619_));
 sky130_fd_sc_hs__nand3_4 _6672_ (.A(_1569_),
    .B(_1571_),
    .C(_1619_),
    .Y(_1620_));
 sky130_fd_sc_hs__and3_1 _6673_ (.A(_3894_),
    .B(_3900_),
    .C(_3887_),
    .X(_1621_));
 sky130_fd_sc_hs__a21oi_4 _6674_ (.A1(_3900_),
    .A2(_3893_),
    .B1(_1621_),
    .Y(_1622_));
 sky130_fd_sc_hs__nor4b_1 _6675_ (.A(_3899_),
    .B(_1084_),
    .C(_1143_),
    .D_N(_3906_),
    .Y(_1623_));
 sky130_fd_sc_hs__a2111oi_2 _6676_ (.A1(_1620_),
    .A2(_1622_),
    .B1(_3906_),
    .C1(_1084_),
    .D1(_1143_),
    .Y(_1624_));
 sky130_fd_sc_hs__a31oi_1 _6677_ (.A1(_1620_),
    .A2(_1622_),
    .A3(_1623_),
    .B1(_1624_),
    .Y(_1625_));
 sky130_fd_sc_hs__nand4b_1 _6678_ (.A_N(_3906_),
    .B(_3899_),
    .C(_1119_),
    .D(_1089_),
    .Y(_1626_));
 sky130_fd_sc_hs__o311ai_2 _6679_ (.A1(_1085_),
    .A2(_1089_),
    .A3(_1318_),
    .B1(_1625_),
    .C1(_1626_),
    .Y(_1627_));
 sky130_fd_sc_hs__a21o_1 _6680_ (.A1(_1606_),
    .A2(_1618_),
    .B1(_1627_),
    .X(net314));
 sky130_fd_sc_hs__a211oi_4 _6681_ (.A1(_0938_),
    .A2(_0975_),
    .B1(_1129_),
    .C1(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[30] ),
    .Y(_1628_));
 sky130_fd_sc_hs__and2_1 _6682_ (.A(_0567_),
    .B(_0932_),
    .X(_1629_));
 sky130_fd_sc_hs__a211oi_2 _6683_ (.A1(net214),
    .A2(_0959_),
    .B1(_1629_),
    .C1(_1210_),
    .Y(_1630_));
 sky130_fd_sc_hs__nor3_1 _6684_ (.A(_3893_),
    .B(_3899_),
    .C(_3905_),
    .Y(_1631_));
 sky130_fd_sc_hs__or2_1 _6685_ (.A(_3906_),
    .B(_3905_),
    .X(_1632_));
 sky130_fd_sc_hs__o31ai_1 _6686_ (.A1(_3900_),
    .A2(_3899_),
    .A3(_3905_),
    .B1(_1632_),
    .Y(_1633_));
 sky130_fd_sc_hs__a31oi_2 _6687_ (.A1(_1589_),
    .A2(_1593_),
    .A3(_1631_),
    .B1(_1633_),
    .Y(_1634_));
 sky130_fd_sc_hs__xnor2_1 _6688_ (.A(_3912_),
    .B(_1634_),
    .Y(_1635_));
 sky130_fd_sc_hs__nand2_1 _6689_ (.A(_1178_),
    .B(_1338_),
    .Y(_1636_));
 sky130_fd_sc_hs__o21ai_2 _6690_ (.A1(_1178_),
    .A2(_1635_),
    .B1(_1636_),
    .Y(_1637_));
 sky130_fd_sc_hs__nand2_8 _6691_ (.A(_1320_),
    .B(_1637_),
    .Y(_1638_));
 sky130_fd_sc_hs__nor2_1 _6692_ (.A(_0567_),
    .B(_1134_),
    .Y(_1639_));
 sky130_fd_sc_hs__nor3_4 _6693_ (.A(_0195_),
    .B(_0196_),
    .C(_1192_),
    .Y(_1640_));
 sky130_fd_sc_hs__a21oi_4 _6694_ (.A1(net144),
    .A2(_1153_),
    .B1(_1154_),
    .Y(_1641_));
 sky130_fd_sc_hs__o21a_1 _6695_ (.A1(_0391_),
    .A2(_1609_),
    .B1(_1641_),
    .X(_1642_));
 sky130_fd_sc_hs__o21ai_1 _6696_ (.A1(_0567_),
    .A2(_1231_),
    .B1(_1241_),
    .Y(_1643_));
 sky130_fd_sc_hs__o32a_1 _6697_ (.A1(_1521_),
    .A2(_1639_),
    .A3(_1640_),
    .B1(_1642_),
    .B2(_1643_),
    .X(_1644_));
 sky130_fd_sc_hs__o311ai_2 _6698_ (.A1(_1082_),
    .A2(_1628_),
    .A3(_1630_),
    .B1(_1638_),
    .C1(_1644_),
    .Y(net315));
 sky130_fd_sc_hs__a21o_1 _6699_ (.A1(net214),
    .A2(_0959_),
    .B1(_1629_),
    .X(_1645_));
 sky130_fd_sc_hs__nor2_2 _6700_ (.A(_1085_),
    .B(_1146_),
    .Y(_1646_));
 sky130_fd_sc_hs__nor3_4 _6701_ (.A(_3899_),
    .B(_3905_),
    .C(_3911_),
    .Y(_1647_));
 sky130_fd_sc_hs__a21oi_2 _6702_ (.A1(_3912_),
    .A2(_1632_),
    .B1(_3911_),
    .Y(_1648_));
 sky130_fd_sc_hs__a31oi_4 _6703_ (.A1(_1620_),
    .A2(_1622_),
    .A3(_1647_),
    .B1(_1648_),
    .Y(_1649_));
 sky130_fd_sc_hs__xnor2_4 _6704_ (.A(_3918_),
    .B(_1649_),
    .Y(_1650_));
 sky130_fd_sc_hs__o2bb2ai_4 _6705_ (.A1_N(_1359_),
    .A2_N(_1646_),
    .B1(_1650_),
    .B2(_1378_),
    .Y(_1651_));
 sky130_fd_sc_hs__nand4_1 _6706_ (.A(_0386_),
    .B(_0382_),
    .C(net215),
    .D(_1079_),
    .Y(_1652_));
 sky130_fd_sc_hs__nand2_1 _6707_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[31] ),
    .B(_1229_),
    .Y(_1653_));
 sky130_fd_sc_hs__nand4_1 _6708_ (.A(_0941_),
    .B(_0974_),
    .C(_0962_),
    .D(_1229_),
    .Y(_1654_));
 sky130_fd_sc_hs__mux2_1 _6709_ (.A0(_0382_),
    .A1(net215),
    .S(_1106_),
    .X(_1655_));
 sky130_fd_sc_hs__a221oi_4 _6710_ (.A1(net145),
    .A2(_0122_),
    .B1(_1655_),
    .B2(_0378_),
    .C1(_1111_),
    .Y(_1656_));
 sky130_fd_sc_hs__o21ai_1 _6711_ (.A1(_0382_),
    .A2(_1114_),
    .B1(_1241_),
    .Y(_1657_));
 sky130_fd_sc_hs__a41oi_2 _6712_ (.A1(_1652_),
    .A2(_1653_),
    .A3(_1654_),
    .A4(_1656_),
    .B1(_1657_),
    .Y(_1658_));
 sky130_fd_sc_hs__a311o_4 _6713_ (.A1(_0103_),
    .A2(_1123_),
    .A3(_1645_),
    .B1(_1651_),
    .C1(_1658_),
    .X(net316));
 sky130_fd_sc_hs__nand3_1 _6714_ (.A(_1264_),
    .B(_0382_),
    .C(net215),
    .Y(_1659_));
 sky130_fd_sc_hs__a31oi_1 _6715_ (.A1(_0430_),
    .A2(net114),
    .A3(_1192_),
    .B1(_1132_),
    .Y(_1660_));
 sky130_fd_sc_hs__nor2_1 _6716_ (.A(net114),
    .B(_1231_),
    .Y(_1661_));
 sky130_fd_sc_hs__a21oi_1 _6717_ (.A1(_1659_),
    .A2(_1660_),
    .B1(_1661_),
    .Y(_1662_));
 sky130_fd_sc_hs__a21o_1 _6718_ (.A1(_3912_),
    .A2(_1634_),
    .B1(_3911_),
    .X(_1663_));
 sky130_fd_sc_hs__a21oi_4 _6719_ (.A1(_3918_),
    .A2(_1663_),
    .B1(_3917_),
    .Y(_1664_));
 sky130_fd_sc_hs__xnor2_4 _6720_ (.A(_3926_),
    .B(_1664_),
    .Y(_1665_));
 sky130_fd_sc_hs__nor2_1 _6721_ (.A(_1086_),
    .B(_1178_),
    .Y(_1666_));
 sky130_fd_sc_hs__a22o_4 _6722_ (.A1(_1328_),
    .A2(_1662_),
    .B1(_1665_),
    .B2(_1666_),
    .X(net317));
 sky130_fd_sc_hs__o21ai_4 _6723_ (.A1(_1109_),
    .A2(_1134_),
    .B1(_1231_),
    .Y(_1667_));
 sky130_fd_sc_hs__nand2_1 _6724_ (.A(net115),
    .B(_1667_),
    .Y(_1668_));
 sky130_fd_sc_hs__nand2_1 _6725_ (.A(_0819_),
    .B(_1668_),
    .Y(_1669_));
 sky130_fd_sc_hs__and2_1 _6726_ (.A(_3926_),
    .B(_3917_),
    .X(_1670_));
 sky130_fd_sc_hs__a311oi_4 _6727_ (.A1(_3926_),
    .A2(_3918_),
    .A3(_1649_),
    .B1(_1670_),
    .C1(_3925_),
    .Y(_1671_));
 sky130_fd_sc_hs__xnor2_1 _6728_ (.A(_2703_),
    .B(_2774_),
    .Y(_1672_));
 sky130_fd_sc_hs__a21oi_1 _6729_ (.A1(net115),
    .A2(_0085_),
    .B1(_0524_),
    .Y(_1673_));
 sky130_fd_sc_hs__xnor2_1 _6730_ (.A(_1672_),
    .B(_1673_),
    .Y(_1674_));
 sky130_fd_sc_hs__xnor2_1 _6731_ (.A(_3547_),
    .B(_2972_),
    .Y(_1675_));
 sky130_fd_sc_hs__xnor2_1 _6732_ (.A(_3545_),
    .B(_3213_),
    .Y(_1676_));
 sky130_fd_sc_hs__xnor2_1 _6733_ (.A(_1675_),
    .B(_1676_),
    .Y(_1677_));
 sky130_fd_sc_hs__xnor2_1 _6734_ (.A(_3922_),
    .B(_3561_),
    .Y(_1678_));
 sky130_fd_sc_hs__xnor2_1 _6735_ (.A(_3549_),
    .B(_3484_),
    .Y(_1679_));
 sky130_fd_sc_hs__xnor2_1 _6736_ (.A(_1678_),
    .B(_1679_),
    .Y(_1680_));
 sky130_fd_sc_hs__xnor2_1 _6737_ (.A(_1677_),
    .B(_1680_),
    .Y(_1681_));
 sky130_fd_sc_hs__xnor2_1 _6738_ (.A(_3552_),
    .B(_3554_),
    .Y(_1682_));
 sky130_fd_sc_hs__xnor2_1 _6739_ (.A(_3543_),
    .B(_3564_),
    .Y(_1683_));
 sky130_fd_sc_hs__xnor2_1 _6740_ (.A(_1682_),
    .B(_1683_),
    .Y(_1684_));
 sky130_fd_sc_hs__xnor2_1 _6741_ (.A(_3485_),
    .B(_3920_),
    .Y(_1685_));
 sky130_fd_sc_hs__xnor2_1 _6742_ (.A(_3558_),
    .B(_1685_),
    .Y(_1686_));
 sky130_fd_sc_hs__xnor2_2 _6743_ (.A(_1684_),
    .B(_1686_),
    .Y(_1687_));
 sky130_fd_sc_hs__xnor2_2 _6744_ (.A(_1681_),
    .B(_1687_),
    .Y(_1688_));
 sky130_fd_sc_hs__xnor2_1 _6745_ (.A(_1674_),
    .B(_1688_),
    .Y(_1689_));
 sky130_fd_sc_hs__xnor2_2 _6746_ (.A(_1671_),
    .B(_1689_),
    .Y(_1690_));
 sky130_fd_sc_hs__o2bb2ai_2 _6747_ (.A1_N(_1606_),
    .A2_N(_1669_),
    .B1(_1690_),
    .B2(_1378_),
    .Y(net318));
 sky130_fd_sc_hs__nand2_1 _6748_ (.A(net219),
    .B(_0989_),
    .Y(_1691_));
 sky130_fd_sc_hs__nand2_1 _6749_ (.A(net181),
    .B(_1035_),
    .Y(_1692_));
 sky130_fd_sc_hs__nor2_1 _6750_ (.A(_0090_),
    .B(net116),
    .Y(_1693_));
 sky130_fd_sc_hs__a311oi_4 _6751_ (.A1(_1037_),
    .A2(_1691_),
    .A3(_1692_),
    .B1(_1693_),
    .C1(_0600_),
    .Y(net319));
 sky130_fd_sc_hs__nand2_1 _6752_ (.A(net220),
    .B(_0989_),
    .Y(_1694_));
 sky130_fd_sc_hs__nand2_1 _6753_ (.A(net182),
    .B(_1035_),
    .Y(_1695_));
 sky130_fd_sc_hs__nor2_1 _6754_ (.A(_0090_),
    .B(net117),
    .Y(_1696_));
 sky130_fd_sc_hs__a311oi_4 _6755_ (.A1(_1037_),
    .A2(_1694_),
    .A3(_1695_),
    .B1(_1696_),
    .C1(_0600_),
    .Y(net320));
 sky130_fd_sc_hs__nand2_1 _6756_ (.A(_0814_),
    .B(net118),
    .Y(_1697_));
 sky130_fd_sc_hs__nand2b_1 _6757_ (.A_N(net183),
    .B(_0992_),
    .Y(_1698_));
 sky130_fd_sc_hs__o211ai_2 _6758_ (.A1(net221),
    .A2(_0993_),
    .B1(_1698_),
    .C1(_1037_),
    .Y(_1699_));
 sky130_fd_sc_hs__a21oi_4 _6759_ (.A1(_1697_),
    .A2(_1699_),
    .B1(_0595_),
    .Y(net321));
 sky130_fd_sc_hs__nor2_1 _6760_ (.A(net184),
    .B(_0989_),
    .Y(_1700_));
 sky130_fd_sc_hs__a211oi_4 _6761_ (.A1(_0299_),
    .A2(_0989_),
    .B1(_1700_),
    .C1(_0813_),
    .Y(_1701_));
 sky130_fd_sc_hs__a21oi_4 _6762_ (.A1(_0814_),
    .A2(net119),
    .B1(_1701_),
    .Y(_1702_));
 sky130_fd_sc_hs__nor2_8 _6763_ (.A(_0109_),
    .B(_1702_),
    .Y(net322));
 sky130_fd_sc_hs__a21oi_4 _6764_ (.A1(_0088_),
    .A2(_0812_),
    .B1(_0595_),
    .Y(net323));
 sky130_fd_sc_hs__nor2_2 _6765_ (.A(_0812_),
    .B(_0109_),
    .Y(net324));
 sky130_fd_sc_hs__nor2_1 _6766_ (.A(_0560_),
    .B(_0548_),
    .Y(_1703_));
 sky130_fd_sc_hs__nor4_2 _6767_ (.A(_0195_),
    .B(_0196_),
    .C(_0560_),
    .D(_0549_),
    .Y(_1704_));
 sky130_fd_sc_hs__or2_1 _6768_ (.A(net14),
    .B(net12),
    .X(_1705_));
 sky130_fd_sc_hs__nor2_1 _6769_ (.A(_0296_),
    .B(_0352_),
    .Y(_1706_));
 sky130_fd_sc_hs__a2111oi_4 _6770_ (.A1(_0247_),
    .A2(_0248_),
    .B1(_0404_),
    .C1(_0408_),
    .D1(_0409_),
    .Y(_1707_));
 sky130_fd_sc_hs__nand4bb_2 _6771_ (.A_N(net198),
    .B_N(net203),
    .C(_1706_),
    .D(_1707_),
    .Y(_1708_));
 sky130_fd_sc_hs__o32ai_1 _6772_ (.A1(_0292_),
    .A2(_0294_),
    .A3(_0295_),
    .B1(_0336_),
    .B2(_0147_),
    .Y(_1709_));
 sky130_fd_sc_hs__o2111ai_2 _6773_ (.A1(_0297_),
    .A2(_0298_),
    .B1(_0309_),
    .C1(_0314_),
    .D1(_0317_),
    .Y(_1710_));
 sky130_fd_sc_hs__nor4_2 _6774_ (.A(net220),
    .B(net217),
    .C(_1709_),
    .D(_1710_),
    .Y(_1711_));
 sky130_fd_sc_hs__a2111oi_1 _6775_ (.A1(_0350_),
    .A2(_0351_),
    .B1(net195),
    .C1(net201),
    .D1(net193),
    .Y(_1712_));
 sky130_fd_sc_hs__o211a_1 _6776_ (.A1(_0333_),
    .A2(_0335_),
    .B1(_0341_),
    .C1(_0345_),
    .X(_1713_));
 sky130_fd_sc_hs__and4b_2 _6777_ (.A_N(net16),
    .B(_1711_),
    .C(_1712_),
    .D(_1713_),
    .X(_1714_));
 sky130_fd_sc_hs__nor4_2 _6778_ (.A(net11),
    .B(net199),
    .C(net206),
    .D(net210),
    .Y(_1715_));
 sky130_fd_sc_hs__nand4bb_2 _6779_ (.A_N(net205),
    .B_N(net204),
    .C(_1714_),
    .D(_1715_),
    .Y(_1716_));
 sky130_fd_sc_hs__nor4_4 _6780_ (.A(net209),
    .B(_1705_),
    .C(_1708_),
    .D(_1716_),
    .Y(_1717_));
 sky130_fd_sc_hs__mux2_1 _6781_ (.A0(_1703_),
    .A1(_1704_),
    .S(_1717_),
    .X(_1718_));
 sky130_fd_sc_hs__nor2_2 _6782_ (.A(_0105_),
    .B(_1142_),
    .Y(_1719_));
 sky130_fd_sc_hs__a22o_2 _6783_ (.A1(_0435_),
    .A2(_1142_),
    .B1(_1719_),
    .B2(_3701_),
    .X(_1720_));
 sky130_fd_sc_hs__a22oi_4 _6784_ (.A1(_0105_),
    .A2(_0435_),
    .B1(_1720_),
    .B2(_0104_),
    .Y(_1721_));
 sky130_fd_sc_hs__o32ai_1 _6785_ (.A1(_0118_),
    .A2(_3570_),
    .A3(_0112_),
    .B1(_0537_),
    .B2(_0532_),
    .Y(_1722_));
 sky130_fd_sc_hs__nand2b_1 _6786_ (.A_N(_3574_),
    .B(_1722_),
    .Y(_1723_));
 sky130_fd_sc_hs__nand2b_1 _6787_ (.A_N(_0532_),
    .B(_0118_),
    .Y(_1724_));
 sky130_fd_sc_hs__a21oi_2 _6788_ (.A1(_0537_),
    .A2(_1724_),
    .B1(_0539_),
    .Y(_1725_));
 sky130_fd_sc_hs__a2bb2oi_4 _6789_ (.A1_N(_0536_),
    .A2_N(_0552_),
    .B1(_1723_),
    .B2(_1725_),
    .Y(_1726_));
 sky130_fd_sc_hs__a221o_1 _6790_ (.A1(_0132_),
    .A2(_1721_),
    .B1(_1703_),
    .B2(net214),
    .C1(_1726_),
    .X(_1727_));
 sky130_fd_sc_hs__nor2_1 _6791_ (.A(_3574_),
    .B(_0112_),
    .Y(_1728_));
 sky130_fd_sc_hs__nor2_2 _6792_ (.A(_0532_),
    .B(_1728_),
    .Y(_1729_));
 sky130_fd_sc_hs__nor2_8 _6793_ (.A(net76),
    .B(net77),
    .Y(_1730_));
 sky130_fd_sc_hs__o211ai_4 _6794_ (.A1(_0118_),
    .A2(_1729_),
    .B1(_1730_),
    .C1(_0537_),
    .Y(_1731_));
 sky130_fd_sc_hs__and3b_4 _6795_ (.A_N(_0110_),
    .B(_0114_),
    .C(_3570_),
    .X(_1732_));
 sky130_fd_sc_hs__nand2_8 _6796_ (.A(_1730_),
    .B(_1732_),
    .Y(_1733_));
 sky130_fd_sc_hs__buf_8 _6797_ (.A(_1733_),
    .X(_1734_));
 sky130_fd_sc_hs__nand2b_4 _6798_ (.A_N(_0537_),
    .B(_1730_),
    .Y(_1735_));
 sky130_fd_sc_hs__nor2_1 _6799_ (.A(_0118_),
    .B(_0112_),
    .Y(_1736_));
 sky130_fd_sc_hs__nor3_4 _6800_ (.A(_0532_),
    .B(_1735_),
    .C(_1736_),
    .Y(_1737_));
 sky130_fd_sc_hs__a21oi_2 _6801_ (.A1(_0532_),
    .A2(_0112_),
    .B1(_3570_),
    .Y(_1738_));
 sky130_fd_sc_hs__a21oi_4 _6802_ (.A1(_0554_),
    .A2(_1738_),
    .B1(_1735_),
    .Y(_1739_));
 sky130_fd_sc_hs__or2_4 _6803_ (.A(net76),
    .B(net77),
    .X(_1740_));
 sky130_fd_sc_hs__nor2_1 _6804_ (.A(_0537_),
    .B(_1740_),
    .Y(_1741_));
 sky130_fd_sc_hs__o211ai_4 _6805_ (.A1(_3574_),
    .A2(_0118_),
    .B1(_1741_),
    .C1(_0532_),
    .Y(_1742_));
 sky130_fd_sc_hs__nor3b_1 _6806_ (.A(_1737_),
    .B(_1739_),
    .C_N(_1742_),
    .Y(_1743_));
 sky130_fd_sc_hs__a41o_4 _6807_ (.A1(_1726_),
    .A2(_1731_),
    .A3(_1734_),
    .A4(_1743_),
    .B1(_0132_),
    .X(_1744_));
 sky130_fd_sc_hs__nand3b_2 _6808_ (.A_N(_0110_),
    .B(_0114_),
    .C(_3570_),
    .Y(_1745_));
 sky130_fd_sc_hs__nor2_8 _6809_ (.A(_1740_),
    .B(_1745_),
    .Y(_1746_));
 sky130_fd_sc_hs__buf_8 _6810_ (.A(_1746_),
    .X(_1747_));
 sky130_fd_sc_hs__clkbuf_8 _6811_ (.A(_1747_),
    .X(_1748_));
 sky130_fd_sc_hs__a31oi_4 _6812_ (.A1(_3948_),
    .A2(_3954_),
    .A3(_3935_),
    .B1(net1),
    .Y(_1749_));
 sky130_fd_sc_hs__xnor2_4 _6813_ (.A(_3960_),
    .B(_1749_),
    .Y(_1750_));
 sky130_fd_sc_hs__buf_8 _6814_ (.A(_1750_),
    .X(_1751_));
 sky130_fd_sc_hs__nand3_4 _6815_ (.A(net2),
    .B(_1730_),
    .C(_1732_),
    .Y(_1752_));
 sky130_fd_sc_hs__o21ai_4 _6816_ (.A1(_1740_),
    .A2(_1745_),
    .B1(net34),
    .Y(_1753_));
 sky130_fd_sc_hs__and2_2 _6817_ (.A(_1752_),
    .B(_1753_),
    .X(_1754_));
 sky130_fd_sc_hs__a31oi_4 _6818_ (.A1(_0562_),
    .A2(_3934_),
    .A3(_3948_),
    .B1(net1),
    .Y(_1755_));
 sky130_fd_sc_hs__xnor2_4 _6819_ (.A(net67),
    .B(_1755_),
    .Y(_1756_));
 sky130_fd_sc_hs__mux2i_4 _6820_ (.A0(_3936_),
    .A1(net53),
    .S(net1),
    .Y(_1757_));
 sky130_fd_sc_hs__clkbuf_16 _6821_ (.A(_1757_),
    .X(_1758_));
 sky130_fd_sc_hs__nor2_8 _6822_ (.A(net1),
    .B(_3935_),
    .Y(_1759_));
 sky130_fd_sc_hs__xnor2_4 _6823_ (.A(net64),
    .B(_1759_),
    .Y(_1760_));
 sky130_fd_sc_hs__nand3_4 _6824_ (.A(_1756_),
    .B(_1758_),
    .C(_1760_),
    .Y(_1761_));
 sky130_fd_sc_hs__nand3_4 _6825_ (.A(_0118_),
    .B(_0545_),
    .C(_1730_),
    .Y(_1762_));
 sky130_fd_sc_hs__o21ai_1 _6826_ (.A1(_0596_),
    .A2(_1761_),
    .B1(_1762_),
    .Y(_1763_));
 sky130_fd_sc_hs__nand2b_4 _6827_ (.A_N(_1754_),
    .B(_1763_),
    .Y(_1764_));
 sky130_fd_sc_hs__a21oi_4 _6828_ (.A1(_1752_),
    .A2(_1753_),
    .B1(_1762_),
    .Y(_1765_));
 sky130_fd_sc_hs__nand2_2 _6829_ (.A(_1750_),
    .B(_1765_),
    .Y(_1766_));
 sky130_fd_sc_hs__o21ai_4 _6830_ (.A1(_1751_),
    .A2(_1764_),
    .B1(_1766_),
    .Y(_1767_));
 sky130_fd_sc_hs__buf_8 _6831_ (.A(_1742_),
    .X(_1768_));
 sky130_fd_sc_hs__nand2_1 _6832_ (.A(_0532_),
    .B(_3570_),
    .Y(_1769_));
 sky130_fd_sc_hs__a21oi_4 _6833_ (.A1(_0554_),
    .A2(_1769_),
    .B1(_1735_),
    .Y(_1770_));
 sky130_fd_sc_hs__clkbuf_4 _6834_ (.A(_1770_),
    .X(_1771_));
 sky130_fd_sc_hs__clkbuf_4 _6835_ (.A(_1771_),
    .X(_1772_));
 sky130_fd_sc_hs__clkbuf_4 _6836_ (.A(_1739_),
    .X(_1773_));
 sky130_fd_sc_hs__o21ai_1 _6837_ (.A1(_3939_),
    .A2(_1772_),
    .B1(_1773_),
    .Y(_1774_));
 sky130_fd_sc_hs__clkbuf_4 _6838_ (.A(_1771_),
    .X(_1775_));
 sky130_fd_sc_hs__or2_2 _6839_ (.A(_1742_),
    .B(_1770_),
    .X(_1776_));
 sky130_fd_sc_hs__buf_4 _6840_ (.A(_1776_),
    .X(_1777_));
 sky130_fd_sc_hs__o2bb2ai_1 _6841_ (.A1_N(_3938_),
    .A2_N(_1775_),
    .B1(_1777_),
    .B2(_3940_),
    .Y(_1778_));
 sky130_fd_sc_hs__a21oi_1 _6842_ (.A1(_1768_),
    .A2(_1774_),
    .B1(_1778_),
    .Y(_1779_));
 sky130_fd_sc_hs__nand2_1 _6843_ (.A(net191),
    .B(_1737_),
    .Y(_1780_));
 sky130_fd_sc_hs__nand2_1 _6844_ (.A(_1721_),
    .B(_1780_),
    .Y(_1781_));
 sky130_fd_sc_hs__a211oi_1 _6845_ (.A1(_1748_),
    .A2(_1767_),
    .B1(_1779_),
    .C1(_1781_),
    .Y(_1782_));
 sky130_fd_sc_hs__mux4_4 _6846_ (.A0(net38),
    .A1(net39),
    .A2(net27),
    .A3(net26),
    .S0(_3933_),
    .S1(_1734_),
    .X(_1783_));
 sky130_fd_sc_hs__buf_8 _6847_ (.A(_1733_),
    .X(_1784_));
 sky130_fd_sc_hs__mux4_4 _6848_ (.A0(net32),
    .A1(net35),
    .A2(net31),
    .A3(net30),
    .S0(_3933_),
    .S1(_1784_),
    .X(_1785_));
 sky130_fd_sc_hs__xnor2_4 _6849_ (.A(_3948_),
    .B(_1759_),
    .Y(_1786_));
 sky130_fd_sc_hs__buf_16 _6850_ (.A(_1786_),
    .X(_1787_));
 sky130_fd_sc_hs__mux2i_4 _6851_ (.A0(_1783_),
    .A1(_1785_),
    .S(_1787_),
    .Y(_1788_));
 sky130_fd_sc_hs__mux4_4 _6852_ (.A0(net36),
    .A1(net37),
    .A2(net29),
    .A3(net28),
    .S0(_3933_),
    .S1(_1734_),
    .X(_1789_));
 sky130_fd_sc_hs__mux4_4 _6853_ (.A0(net34),
    .A1(net2),
    .A2(net33),
    .A3(net21),
    .S0(_1746_),
    .S1(_3933_),
    .X(_1790_));
 sky130_fd_sc_hs__mux2i_4 _6854_ (.A0(_1789_),
    .A1(_1790_),
    .S(_1787_),
    .Y(_1791_));
 sky130_fd_sc_hs__mux2_1 _6855_ (.A0(_3936_),
    .A1(net53),
    .S(net1),
    .X(_1792_));
 sky130_fd_sc_hs__buf_8 _6856_ (.A(_1792_),
    .X(_1793_));
 sky130_fd_sc_hs__clkbuf_16 _6857_ (.A(_1793_),
    .X(_1794_));
 sky130_fd_sc_hs__mux2i_4 _6858_ (.A0(_1788_),
    .A1(_1791_),
    .S(_1794_),
    .Y(_1795_));
 sky130_fd_sc_hs__mux4_4 _6859_ (.A0(net5),
    .A1(net6),
    .A2(net20),
    .A3(net19),
    .S0(_0563_),
    .S1(_1784_),
    .X(_1796_));
 sky130_fd_sc_hs__mux4_4 _6860_ (.A0(net40),
    .A1(net41),
    .A2(net25),
    .A3(net24),
    .S0(_0563_),
    .S1(_1784_),
    .X(_1797_));
 sky130_fd_sc_hs__mux2i_4 _6861_ (.A0(_1796_),
    .A1(_1797_),
    .S(_1786_),
    .Y(_1798_));
 sky130_fd_sc_hs__mux4_4 _6862_ (.A0(net7),
    .A1(net8),
    .A2(net18),
    .A3(net17),
    .S0(_0563_),
    .S1(_1784_),
    .X(_1799_));
 sky130_fd_sc_hs__mux4_4 _6863_ (.A0(net3),
    .A1(net4),
    .A2(net23),
    .A3(net22),
    .S0(_0563_),
    .S1(_1784_),
    .X(_1800_));
 sky130_fd_sc_hs__mux2i_4 _6864_ (.A0(_1799_),
    .A1(_1800_),
    .S(_1786_),
    .Y(_1801_));
 sky130_fd_sc_hs__mux2i_4 _6865_ (.A0(_1798_),
    .A1(_1801_),
    .S(_1758_),
    .Y(_1802_));
 sky130_fd_sc_hs__buf_8 _6866_ (.A(_1756_),
    .X(_1803_));
 sky130_fd_sc_hs__mux2i_4 _6867_ (.A0(_1795_),
    .A1(_1802_),
    .S(_1803_),
    .Y(_1804_));
 sky130_fd_sc_hs__buf_8 _6868_ (.A(_1756_),
    .X(_1805_));
 sky130_fd_sc_hs__buf_8 _6869_ (.A(_1786_),
    .X(_1806_));
 sky130_fd_sc_hs__clkbuf_16 _6870_ (.A(_0561_),
    .X(_1807_));
 sky130_fd_sc_hs__buf_8 _6871_ (.A(_1746_),
    .X(_1808_));
 sky130_fd_sc_hs__mux4_4 _6872_ (.A0(net36),
    .A1(net37),
    .A2(net29),
    .A3(net28),
    .S0(_1807_),
    .S1(_1808_),
    .X(_1809_));
 sky130_fd_sc_hs__mux4_4 _6873_ (.A0(net38),
    .A1(net39),
    .A2(net27),
    .A3(net26),
    .S0(_0596_),
    .S1(_1747_),
    .X(_1810_));
 sky130_fd_sc_hs__mux2i_4 _6874_ (.A0(_1809_),
    .A1(_1810_),
    .S(_1794_),
    .Y(_1811_));
 sky130_fd_sc_hs__nand2_1 _6875_ (.A(_1806_),
    .B(_1811_),
    .Y(_1812_));
 sky130_fd_sc_hs__a21oi_1 _6876_ (.A1(_1730_),
    .A2(_1732_),
    .B1(_3953_),
    .Y(_1813_));
 sky130_fd_sc_hs__a21oi_2 _6877_ (.A1(net30),
    .A2(_1808_),
    .B1(_1813_),
    .Y(_1814_));
 sky130_fd_sc_hs__a21oi_2 _6878_ (.A1(_1730_),
    .A2(_1732_),
    .B1(_3947_),
    .Y(_1815_));
 sky130_fd_sc_hs__a21oi_4 _6879_ (.A1(net31),
    .A2(_1808_),
    .B1(_1815_),
    .Y(_1816_));
 sky130_fd_sc_hs__mux2i_4 _6880_ (.A0(_1814_),
    .A1(_1816_),
    .S(_3933_),
    .Y(_1817_));
 sky130_fd_sc_hs__a21oi_1 _6881_ (.A1(_1730_),
    .A2(_1732_),
    .B1(_3942_),
    .Y(_1818_));
 sky130_fd_sc_hs__a21oi_1 _6882_ (.A1(net33),
    .A2(_1808_),
    .B1(_1818_),
    .Y(_1819_));
 sky130_fd_sc_hs__nor2_1 _6883_ (.A(_3927_),
    .B(_1784_),
    .Y(_1820_));
 sky130_fd_sc_hs__a211oi_1 _6884_ (.A1(net2),
    .A2(_1784_),
    .B1(_1820_),
    .C1(_0596_),
    .Y(_1821_));
 sky130_fd_sc_hs__clkbuf_16 _6885_ (.A(_1793_),
    .X(_1822_));
 sky130_fd_sc_hs__a211oi_1 _6886_ (.A1(_0596_),
    .A2(_1819_),
    .B1(_1821_),
    .C1(_1822_),
    .Y(_1823_));
 sky130_fd_sc_hs__a211o_2 _6887_ (.A1(_1794_),
    .A2(_1817_),
    .B1(_1823_),
    .C1(_1806_),
    .X(_1824_));
 sky130_fd_sc_hs__mux4_4 _6888_ (.A0(net40),
    .A1(net41),
    .A2(net25),
    .A3(net24),
    .S0(_1807_),
    .S1(_1746_),
    .X(_1825_));
 sky130_fd_sc_hs__mux4_4 _6889_ (.A0(net3),
    .A1(net4),
    .A2(net23),
    .A3(net22),
    .S0(_1807_),
    .S1(_1808_),
    .X(_1826_));
 sky130_fd_sc_hs__mux2i_4 _6890_ (.A0(_1825_),
    .A1(_1826_),
    .S(_1793_),
    .Y(_1827_));
 sky130_fd_sc_hs__mux4_4 _6891_ (.A0(net5),
    .A1(net6),
    .A2(net20),
    .A3(net19),
    .S0(_1807_),
    .S1(_1808_),
    .X(_1828_));
 sky130_fd_sc_hs__mux4_4 _6892_ (.A0(net7),
    .A1(net8),
    .A2(net18),
    .A3(net17),
    .S0(_1807_),
    .S1(_1808_),
    .X(_1829_));
 sky130_fd_sc_hs__mux2i_4 _6893_ (.A0(_1828_),
    .A1(_1829_),
    .S(_1793_),
    .Y(_1830_));
 sky130_fd_sc_hs__mux2i_4 _6894_ (.A0(_1827_),
    .A1(_1830_),
    .S(_1787_),
    .Y(_1831_));
 sky130_fd_sc_hs__nor2b_1 _6895_ (.A(_1756_),
    .B_N(_1831_),
    .Y(_1832_));
 sky130_fd_sc_hs__a311oi_4 _6896_ (.A1(_1805_),
    .A2(_1812_),
    .A3(_1824_),
    .B1(_1832_),
    .C1(_1750_),
    .Y(_1833_));
 sky130_fd_sc_hs__a21oi_4 _6897_ (.A1(_1751_),
    .A2(_1804_),
    .B1(_1833_),
    .Y(_1834_));
 sky130_fd_sc_hs__nor2_8 _6898_ (.A(_1731_),
    .B(_1732_),
    .Y(_1835_));
 sky130_fd_sc_hs__buf_8 _6899_ (.A(_1835_),
    .X(_1836_));
 sky130_fd_sc_hs__nand2_1 _6900_ (.A(_1834_),
    .B(_1836_),
    .Y(_1837_));
 sky130_fd_sc_hs__a22o_2 _6901_ (.A1(_1721_),
    .A2(_1744_),
    .B1(_1782_),
    .B2(_1837_),
    .X(_1838_));
 sky130_fd_sc_hs__o21ai_4 _6902_ (.A1(_1718_),
    .A2(_1727_),
    .B1(_1838_),
    .Y(net325));
 sky130_fd_sc_hs__clkbuf_16 _6903_ (.A(_1744_),
    .X(_1839_));
 sky130_fd_sc_hs__buf_8 _6904_ (.A(_1737_),
    .X(_1840_));
 sky130_fd_sc_hs__clkbuf_8 _6905_ (.A(_1747_),
    .X(_1841_));
 sky130_fd_sc_hs__xnor2_4 _6906_ (.A(net68),
    .B(_1749_),
    .Y(_1842_));
 sky130_fd_sc_hs__clkbuf_16 _6907_ (.A(_1842_),
    .X(_1843_));
 sky130_fd_sc_hs__clkbuf_16 _6908_ (.A(_1756_),
    .X(_1844_));
 sky130_fd_sc_hs__mux4_4 _6909_ (.A0(net37),
    .A1(net38),
    .A2(net28),
    .A3(net27),
    .S0(_0563_),
    .S1(_1784_),
    .X(_1845_));
 sky130_fd_sc_hs__mux4_4 _6910_ (.A0(net35),
    .A1(net36),
    .A2(net30),
    .A3(net29),
    .S0(_3933_),
    .S1(_1734_),
    .X(_1846_));
 sky130_fd_sc_hs__mux2i_4 _6911_ (.A0(_1845_),
    .A1(_1846_),
    .S(_1822_),
    .Y(_1847_));
 sky130_fd_sc_hs__mux4_4 _6912_ (.A0(net41),
    .A1(net3),
    .A2(net24),
    .A3(net23),
    .S0(_0563_),
    .S1(_1733_),
    .X(_1848_));
 sky130_fd_sc_hs__mux4_4 _6913_ (.A0(net39),
    .A1(net40),
    .A2(net26),
    .A3(net25),
    .S0(_0563_),
    .S1(_1733_),
    .X(_1849_));
 sky130_fd_sc_hs__mux2i_4 _6914_ (.A0(_1848_),
    .A1(_1849_),
    .S(_1822_),
    .Y(_1850_));
 sky130_fd_sc_hs__clkbuf_16 _6915_ (.A(_1760_),
    .X(_1851_));
 sky130_fd_sc_hs__mux2i_4 _6916_ (.A0(_1847_),
    .A1(_1850_),
    .S(_1851_),
    .Y(_1852_));
 sky130_fd_sc_hs__mux4_4 _6917_ (.A0(net21),
    .A1(net32),
    .A2(net33),
    .A3(net31),
    .S0(_3933_),
    .S1(_1784_),
    .X(_1853_));
 sky130_fd_sc_hs__a22oi_4 _6918_ (.A1(_1752_),
    .A2(_1753_),
    .B1(_1762_),
    .B2(_0596_),
    .Y(_1854_));
 sky130_fd_sc_hs__mux2i_4 _6919_ (.A0(_1853_),
    .A1(_1854_),
    .S(_1793_),
    .Y(_1855_));
 sky130_fd_sc_hs__nor2_4 _6920_ (.A(_1765_),
    .B(_1851_),
    .Y(_1856_));
 sky130_fd_sc_hs__a211oi_4 _6921_ (.A1(_1851_),
    .A2(_1855_),
    .B1(_1856_),
    .C1(_1803_),
    .Y(_1857_));
 sky130_fd_sc_hs__a21oi_4 _6922_ (.A1(_1844_),
    .A2(_1852_),
    .B1(_1857_),
    .Y(_1858_));
 sky130_fd_sc_hs__nor2_4 _6923_ (.A(_1842_),
    .B(_1765_),
    .Y(_1859_));
 sky130_fd_sc_hs__buf_8 _6924_ (.A(_1859_),
    .X(_1860_));
 sky130_fd_sc_hs__a21oi_4 _6925_ (.A1(_1843_),
    .A2(_1858_),
    .B1(_1860_),
    .Y(_1861_));
 sky130_fd_sc_hs__buf_8 _6926_ (.A(_1756_),
    .X(_1862_));
 sky130_fd_sc_hs__mux2i_4 _6927_ (.A0(_1765_),
    .A1(_1785_),
    .S(_1760_),
    .Y(_1863_));
 sky130_fd_sc_hs__mux2i_4 _6928_ (.A0(_1791_),
    .A1(_1863_),
    .S(_1794_),
    .Y(_1864_));
 sky130_fd_sc_hs__nor3_4 _6929_ (.A(_1754_),
    .B(_1762_),
    .C(_1756_),
    .Y(_1865_));
 sky130_fd_sc_hs__a21oi_4 _6930_ (.A1(_1862_),
    .A2(_1864_),
    .B1(_1865_),
    .Y(_1866_));
 sky130_fd_sc_hs__mux2i_4 _6931_ (.A0(_1800_),
    .A1(_1783_),
    .S(_1787_),
    .Y(_1867_));
 sky130_fd_sc_hs__mux2i_4 _6932_ (.A0(_1798_),
    .A1(_1867_),
    .S(_1794_),
    .Y(_1868_));
 sky130_fd_sc_hs__mux2i_4 _6933_ (.A0(_1826_),
    .A1(_1828_),
    .S(_1793_),
    .Y(_1869_));
 sky130_fd_sc_hs__mux2i_4 _6934_ (.A0(_1799_),
    .A1(_1829_),
    .S(_1757_),
    .Y(_1870_));
 sky130_fd_sc_hs__mux2i_4 _6935_ (.A0(_1869_),
    .A1(_1870_),
    .S(_1787_),
    .Y(_1871_));
 sky130_fd_sc_hs__mux2i_4 _6936_ (.A0(_1868_),
    .A1(_1871_),
    .S(_1862_),
    .Y(_1872_));
 sky130_fd_sc_hs__mux2i_4 _6937_ (.A0(_1866_),
    .A1(_1872_),
    .S(_1843_),
    .Y(_1873_));
 sky130_fd_sc_hs__clkbuf_8 _6938_ (.A(_1835_),
    .X(_1874_));
 sky130_fd_sc_hs__clkbuf_16 _6939_ (.A(_1742_),
    .X(_1875_));
 sky130_fd_sc_hs__buf_4 _6940_ (.A(_1739_),
    .X(_1876_));
 sky130_fd_sc_hs__o21ai_1 _6941_ (.A1(_3998_),
    .A2(_1775_),
    .B1(_1876_),
    .Y(_1877_));
 sky130_fd_sc_hs__o2bb2ai_1 _6942_ (.A1_N(_3997_),
    .A2_N(_1775_),
    .B1(_1777_),
    .B2(_3999_),
    .Y(_1878_));
 sky130_fd_sc_hs__a21oi_2 _6943_ (.A1(_1875_),
    .A2(_1877_),
    .B1(_1878_),
    .Y(_1879_));
 sky130_fd_sc_hs__a221o_1 _6944_ (.A1(_1841_),
    .A2(_1861_),
    .B1(_1873_),
    .B2(_1874_),
    .C1(_1879_),
    .X(_1880_));
 sky130_fd_sc_hs__a21oi_2 _6945_ (.A1(net192),
    .A2(_1840_),
    .B1(_1880_),
    .Y(_1881_));
 sky130_fd_sc_hs__a21oi_1 _6946_ (.A1(_1242_),
    .A2(_0580_),
    .B1(_1276_),
    .Y(_1882_));
 sky130_fd_sc_hs__o21ai_4 _6947_ (.A1(_1839_),
    .A2(_1881_),
    .B1(_1882_),
    .Y(net326));
 sky130_fd_sc_hs__mux2i_4 _6948_ (.A0(_1797_),
    .A1(_1789_),
    .S(_1787_),
    .Y(_1883_));
 sky130_fd_sc_hs__mux2i_4 _6949_ (.A0(_1867_),
    .A1(_1883_),
    .S(_1794_),
    .Y(_1884_));
 sky130_fd_sc_hs__buf_8 _6950_ (.A(_1760_),
    .X(_1885_));
 sky130_fd_sc_hs__mux2i_4 _6951_ (.A0(_1785_),
    .A1(_1790_),
    .S(_1822_),
    .Y(_1886_));
 sky130_fd_sc_hs__a211oi_4 _6952_ (.A1(_1885_),
    .A2(_1886_),
    .B1(_1856_),
    .C1(_1803_),
    .Y(_1887_));
 sky130_fd_sc_hs__a21oi_4 _6953_ (.A1(_1862_),
    .A2(_1884_),
    .B1(_1887_),
    .Y(_1888_));
 sky130_fd_sc_hs__a21oi_4 _6954_ (.A1(_1843_),
    .A2(_1888_),
    .B1(_1860_),
    .Y(_1889_));
 sky130_fd_sc_hs__clkbuf_16 _6955_ (.A(_1842_),
    .X(_1890_));
 sky130_fd_sc_hs__mux4_4 _6956_ (.A0(net4),
    .A1(net5),
    .A2(net22),
    .A3(net20),
    .S0(_0563_),
    .S1(_1733_),
    .X(_1891_));
 sky130_fd_sc_hs__mux4_4 _6957_ (.A0(_1845_),
    .A1(_1848_),
    .A2(_1849_),
    .A3(_1891_),
    .S0(_1760_),
    .S1(_1757_),
    .X(_1892_));
 sky130_fd_sc_hs__inv_1 _6958_ (.A(_1892_),
    .Y(_1893_));
 sky130_fd_sc_hs__mux4_4 _6959_ (.A0(net6),
    .A1(net7),
    .A2(net19),
    .A3(net18),
    .S0(_0563_),
    .S1(_1784_),
    .X(_1894_));
 sky130_fd_sc_hs__nor2_1 _6960_ (.A(_1757_),
    .B(_1894_),
    .Y(_1895_));
 sky130_fd_sc_hs__xnor2_4 _6961_ (.A(_3933_),
    .B(_1746_),
    .Y(_1896_));
 sky130_fd_sc_hs__mux2i_4 _6962_ (.A0(_4025_),
    .A1(_4031_),
    .S(_1896_),
    .Y(_1897_));
 sky130_fd_sc_hs__nor2_1 _6963_ (.A(_1822_),
    .B(_1897_),
    .Y(_1898_));
 sky130_fd_sc_hs__mux4_4 _6964_ (.A0(net4),
    .A1(net5),
    .A2(net22),
    .A3(net20),
    .S0(_1807_),
    .S1(_1746_),
    .X(_1899_));
 sky130_fd_sc_hs__mux4_4 _6965_ (.A0(net6),
    .A1(net7),
    .A2(net19),
    .A3(net18),
    .S0(_1807_),
    .S1(_1746_),
    .X(_1900_));
 sky130_fd_sc_hs__mux2_1 _6966_ (.A0(_1899_),
    .A1(_1900_),
    .S(_1793_),
    .X(_1901_));
 sky130_fd_sc_hs__nand2_1 _6967_ (.A(_1851_),
    .B(_1901_),
    .Y(_1902_));
 sky130_fd_sc_hs__o31a_1 _6968_ (.A1(_1760_),
    .A2(_1895_),
    .A3(_1898_),
    .B1(_1902_),
    .X(_1903_));
 sky130_fd_sc_hs__mux2_1 _6969_ (.A0(_1893_),
    .A1(_1903_),
    .S(_1805_),
    .X(_1904_));
 sky130_fd_sc_hs__o21ai_1 _6970_ (.A1(_0596_),
    .A2(_1793_),
    .B1(_1762_),
    .Y(_1905_));
 sky130_fd_sc_hs__nand2_1 _6971_ (.A(_1787_),
    .B(_1905_),
    .Y(_1906_));
 sky130_fd_sc_hs__mux2i_4 _6972_ (.A0(_1846_),
    .A1(_1853_),
    .S(_1822_),
    .Y(_1907_));
 sky130_fd_sc_hs__o22ai_4 _6973_ (.A1(_1754_),
    .A2(_1906_),
    .B1(_1907_),
    .B2(_1806_),
    .Y(_1908_));
 sky130_fd_sc_hs__a211oi_4 _6974_ (.A1(_1862_),
    .A2(_1908_),
    .B1(_1865_),
    .C1(_1842_),
    .Y(_1909_));
 sky130_fd_sc_hs__a21oi_4 _6975_ (.A1(_1890_),
    .A2(_1904_),
    .B1(_1909_),
    .Y(_1910_));
 sky130_fd_sc_hs__o21ai_1 _6976_ (.A1(_4004_),
    .A2(_1775_),
    .B1(_1876_),
    .Y(_1911_));
 sky130_fd_sc_hs__clkbuf_4 _6977_ (.A(_1771_),
    .X(_1912_));
 sky130_fd_sc_hs__o2bb2ai_1 _6978_ (.A1_N(_4003_),
    .A2_N(_1912_),
    .B1(_1777_),
    .B2(_4005_),
    .Y(_1913_));
 sky130_fd_sc_hs__a21oi_4 _6979_ (.A1(_1875_),
    .A2(_1911_),
    .B1(_1913_),
    .Y(_1914_));
 sky130_fd_sc_hs__a221o_1 _6980_ (.A1(_1841_),
    .A2(_1889_),
    .B1(_1910_),
    .B2(_1874_),
    .C1(_1914_),
    .X(_1915_));
 sky130_fd_sc_hs__a21oi_2 _6981_ (.A1(net365),
    .A2(_1840_),
    .B1(_1915_),
    .Y(_1916_));
 sky130_fd_sc_hs__a21oi_1 _6982_ (.A1(_1242_),
    .A2(_0581_),
    .B1(_1284_),
    .Y(_1917_));
 sky130_fd_sc_hs__o21ai_4 _6983_ (.A1(_1839_),
    .A2(_1916_),
    .B1(_1917_),
    .Y(net327));
 sky130_fd_sc_hs__mux2i_4 _6984_ (.A0(_1908_),
    .A1(_1892_),
    .S(_1803_),
    .Y(_1918_));
 sky130_fd_sc_hs__a21oi_2 _6985_ (.A1(_1843_),
    .A2(_1918_),
    .B1(_1859_),
    .Y(_1919_));
 sky130_fd_sc_hs__nand2b_4 _6986_ (.A_N(_1731_),
    .B(_1745_),
    .Y(_1920_));
 sky130_fd_sc_hs__and2_1 _6987_ (.A(_1793_),
    .B(_1796_),
    .X(_1921_));
 sky130_fd_sc_hs__a211oi_4 _6988_ (.A1(_1758_),
    .A2(_1799_),
    .B1(_1921_),
    .C1(_1760_),
    .Y(_1922_));
 sky130_fd_sc_hs__a21oi_4 _6989_ (.A1(_1851_),
    .A2(_1830_),
    .B1(_1922_),
    .Y(_1923_));
 sky130_fd_sc_hs__mux2_1 _6990_ (.A0(_1884_),
    .A1(_1923_),
    .S(_1803_),
    .X(_1924_));
 sky130_fd_sc_hs__a21oi_4 _6991_ (.A1(_1803_),
    .A2(_1851_),
    .B1(_1765_),
    .Y(_1925_));
 sky130_fd_sc_hs__a311oi_4 _6992_ (.A1(_1862_),
    .A2(_1885_),
    .A3(_1886_),
    .B1(_1925_),
    .C1(_1842_),
    .Y(_1926_));
 sky130_fd_sc_hs__a21oi_4 _6993_ (.A1(_1890_),
    .A2(_1924_),
    .B1(_1926_),
    .Y(_1927_));
 sky130_fd_sc_hs__clkbuf_4 _6994_ (.A(_1737_),
    .X(_1928_));
 sky130_fd_sc_hs__o21ai_1 _6995_ (.A1(_4010_),
    .A2(_1772_),
    .B1(_1773_),
    .Y(_1929_));
 sky130_fd_sc_hs__buf_4 _6996_ (.A(_1776_),
    .X(_1930_));
 sky130_fd_sc_hs__o2bb2ai_1 _6997_ (.A1_N(_4009_),
    .A2_N(_1772_),
    .B1(_1930_),
    .B2(_4011_),
    .Y(_1931_));
 sky130_fd_sc_hs__a21oi_2 _6998_ (.A1(_1768_),
    .A2(_1929_),
    .B1(_1931_),
    .Y(_1932_));
 sky130_fd_sc_hs__a21oi_1 _6999_ (.A1(net194),
    .A2(_1928_),
    .B1(_1932_),
    .Y(_1933_));
 sky130_fd_sc_hs__o21ai_1 _7000_ (.A1(_1920_),
    .A2(_1927_),
    .B1(_1933_),
    .Y(_1934_));
 sky130_fd_sc_hs__a21oi_2 _7001_ (.A1(_1748_),
    .A2(_1919_),
    .B1(_1934_),
    .Y(_1935_));
 sky130_fd_sc_hs__a21oi_4 _7002_ (.A1(_1242_),
    .A2(_0582_),
    .B1(_1305_),
    .Y(_1936_));
 sky130_fd_sc_hs__o21ai_4 _7003_ (.A1(_1839_),
    .A2(_1935_),
    .B1(_1936_),
    .Y(net328));
 sky130_fd_sc_hs__clkbuf_16 _7004_ (.A(_1744_),
    .X(_1937_));
 sky130_fd_sc_hs__clkbuf_4 _7005_ (.A(_1771_),
    .X(_1938_));
 sky130_fd_sc_hs__o21ai_1 _7006_ (.A1(_4016_),
    .A2(_1938_),
    .B1(_1773_),
    .Y(_1939_));
 sky130_fd_sc_hs__o2bb2ai_1 _7007_ (.A1_N(_4015_),
    .A2_N(_1938_),
    .B1(_1930_),
    .B2(_4017_),
    .Y(_1940_));
 sky130_fd_sc_hs__a21oi_2 _7008_ (.A1(_1768_),
    .A2(_1939_),
    .B1(_1940_),
    .Y(_1941_));
 sky130_fd_sc_hs__mux2i_4 _7009_ (.A0(_1864_),
    .A1(_1868_),
    .S(_1805_),
    .Y(_1942_));
 sky130_fd_sc_hs__a21oi_4 _7010_ (.A1(_1890_),
    .A2(_1942_),
    .B1(_1860_),
    .Y(_1943_));
 sky130_fd_sc_hs__a31oi_4 _7011_ (.A1(_1844_),
    .A2(_1885_),
    .A3(_1855_),
    .B1(_1925_),
    .Y(_1944_));
 sky130_fd_sc_hs__mux2i_4 _7012_ (.A0(_1900_),
    .A1(_1897_),
    .S(_1794_),
    .Y(_1945_));
 sky130_fd_sc_hs__mux2i_4 _7013_ (.A0(_1894_),
    .A1(_1891_),
    .S(_1822_),
    .Y(_1946_));
 sky130_fd_sc_hs__mux2i_4 _7014_ (.A0(_1945_),
    .A1(_1946_),
    .S(_1806_),
    .Y(_1947_));
 sky130_fd_sc_hs__mux2_1 _7015_ (.A0(_1852_),
    .A1(_1947_),
    .S(_1844_),
    .X(_1948_));
 sky130_fd_sc_hs__mux2i_4 _7016_ (.A0(_1944_),
    .A1(_1948_),
    .S(_1890_),
    .Y(_1949_));
 sky130_fd_sc_hs__o2bb2ai_2 _7017_ (.A1_N(_1748_),
    .A2_N(_1943_),
    .B1(_1949_),
    .B2(_1920_),
    .Y(_1950_));
 sky130_fd_sc_hs__a211oi_4 _7018_ (.A1(net195),
    .A2(_1840_),
    .B1(_1941_),
    .C1(_1950_),
    .Y(_1951_));
 sky130_fd_sc_hs__nand2_1 _7019_ (.A(_1606_),
    .B(_0584_),
    .Y(_1952_));
 sky130_fd_sc_hs__o211ai_4 _7020_ (.A1(_1937_),
    .A2(_1951_),
    .B1(_1952_),
    .C1(_1321_),
    .Y(net329));
 sky130_fd_sc_hs__buf_8 _7021_ (.A(_1737_),
    .X(_1953_));
 sky130_fd_sc_hs__mux2i_4 _7022_ (.A0(_1847_),
    .A1(_1855_),
    .S(_1787_),
    .Y(_1954_));
 sky130_fd_sc_hs__mux2i_4 _7023_ (.A0(_1850_),
    .A1(_1946_),
    .S(_1851_),
    .Y(_1955_));
 sky130_fd_sc_hs__mux2i_4 _7024_ (.A0(_1954_),
    .A1(_1955_),
    .S(_1803_),
    .Y(_1956_));
 sky130_fd_sc_hs__a211oi_4 _7025_ (.A1(_1890_),
    .A2(_1956_),
    .B1(_1860_),
    .C1(_1734_),
    .Y(_1957_));
 sky130_fd_sc_hs__o21ai_1 _7026_ (.A1(_4022_),
    .A2(_1938_),
    .B1(_1773_),
    .Y(_1958_));
 sky130_fd_sc_hs__o2bb2ai_1 _7027_ (.A1_N(_4021_),
    .A2_N(_1938_),
    .B1(_1930_),
    .B2(_4023_),
    .Y(_1959_));
 sky130_fd_sc_hs__a21oi_2 _7028_ (.A1(_1768_),
    .A2(_1958_),
    .B1(_1959_),
    .Y(_1960_));
 sky130_fd_sc_hs__mux2i_4 _7029_ (.A0(_1790_),
    .A1(_1765_),
    .S(_1761_),
    .Y(_1961_));
 sky130_fd_sc_hs__mux2i_4 _7030_ (.A0(_1788_),
    .A1(_1883_),
    .S(_1758_),
    .Y(_1962_));
 sky130_fd_sc_hs__and2_1 _7031_ (.A(_1757_),
    .B(_1796_),
    .X(_1963_));
 sky130_fd_sc_hs__a211oi_4 _7032_ (.A1(_1794_),
    .A2(_1800_),
    .B1(_1963_),
    .C1(_1851_),
    .Y(_1964_));
 sky130_fd_sc_hs__a21oi_4 _7033_ (.A1(_1885_),
    .A2(_1870_),
    .B1(_1964_),
    .Y(_1965_));
 sky130_fd_sc_hs__mux2i_1 _7034_ (.A0(_1962_),
    .A1(_1965_),
    .S(_1844_),
    .Y(_1966_));
 sky130_fd_sc_hs__mux2_2 _7035_ (.A0(_1961_),
    .A1(_1966_),
    .S(_1842_),
    .X(_1967_));
 sky130_fd_sc_hs__nor2_1 _7036_ (.A(_1920_),
    .B(_1967_),
    .Y(_1968_));
 sky130_fd_sc_hs__a2111oi_4 _7037_ (.A1(net196),
    .A2(_1953_),
    .B1(_1957_),
    .C1(_1960_),
    .D1(_1968_),
    .Y(_1969_));
 sky130_fd_sc_hs__a21oi_2 _7038_ (.A1(_1242_),
    .A2(_0585_),
    .B1(_1340_),
    .Y(_1970_));
 sky130_fd_sc_hs__o21ai_4 _7039_ (.A1(_1839_),
    .A2(_1969_),
    .B1(_1970_),
    .Y(net330));
 sky130_fd_sc_hs__mux2i_4 _7040_ (.A0(_1845_),
    .A1(_1853_),
    .S(_1787_),
    .Y(_1971_));
 sky130_fd_sc_hs__mux2i_4 _7041_ (.A0(_1846_),
    .A1(_1849_),
    .S(_1760_),
    .Y(_1972_));
 sky130_fd_sc_hs__mux2i_4 _7042_ (.A0(_1971_),
    .A1(_1972_),
    .S(_1758_),
    .Y(_1973_));
 sky130_fd_sc_hs__mux4_2 _7043_ (.A0(_1848_),
    .A1(_1894_),
    .A2(_1891_),
    .A3(_1897_),
    .S0(_1760_),
    .S1(_1758_),
    .X(_1974_));
 sky130_fd_sc_hs__mux2i_4 _7044_ (.A0(_1973_),
    .A1(_1974_),
    .S(_1805_),
    .Y(_1975_));
 sky130_fd_sc_hs__mux2i_4 _7045_ (.A0(_1764_),
    .A1(_1975_),
    .S(_1842_),
    .Y(_1976_));
 sky130_fd_sc_hs__a22oi_2 _7046_ (.A1(net197),
    .A2(_1928_),
    .B1(_1836_),
    .B2(_1976_),
    .Y(_1977_));
 sky130_fd_sc_hs__a21oi_4 _7047_ (.A1(_1890_),
    .A2(_1804_),
    .B1(_1860_),
    .Y(_1978_));
 sky130_fd_sc_hs__o21ai_1 _7048_ (.A1(_4028_),
    .A2(_1772_),
    .B1(_1773_),
    .Y(_1979_));
 sky130_fd_sc_hs__o2bb2ai_1 _7049_ (.A1_N(_4027_),
    .A2_N(_1772_),
    .B1(_1930_),
    .B2(_4029_),
    .Y(_1980_));
 sky130_fd_sc_hs__a21oi_1 _7050_ (.A1(_1768_),
    .A2(_1979_),
    .B1(_1980_),
    .Y(_1981_));
 sky130_fd_sc_hs__a21oi_2 _7051_ (.A1(_1748_),
    .A2(_1978_),
    .B1(_1981_),
    .Y(_1982_));
 sky130_fd_sc_hs__clkbuf_8 _7052_ (.A(_1744_),
    .X(_1983_));
 sky130_fd_sc_hs__a21oi_4 _7053_ (.A1(_1977_),
    .A2(_1982_),
    .B1(_1983_),
    .Y(_1984_));
 sky130_fd_sc_hs__a21oi_4 _7054_ (.A1(_1242_),
    .A2(net107),
    .B1(_1984_),
    .Y(_1985_));
 sky130_fd_sc_hs__nand2_8 _7055_ (.A(_1362_),
    .B(_1985_),
    .Y(net331));
 sky130_fd_sc_hs__buf_8 _7056_ (.A(_1742_),
    .X(_1986_));
 sky130_fd_sc_hs__clkbuf_4 _7057_ (.A(_1771_),
    .X(_1987_));
 sky130_fd_sc_hs__clkbuf_4 _7058_ (.A(_1739_),
    .X(_1988_));
 sky130_fd_sc_hs__o21ai_1 _7059_ (.A1(_4034_),
    .A2(_1987_),
    .B1(_1988_),
    .Y(_1989_));
 sky130_fd_sc_hs__buf_4 _7060_ (.A(_1776_),
    .X(_1990_));
 sky130_fd_sc_hs__o2bb2ai_1 _7061_ (.A1_N(_4033_),
    .A2_N(_1987_),
    .B1(_1990_),
    .B2(_4035_),
    .Y(_1991_));
 sky130_fd_sc_hs__a21oi_4 _7062_ (.A1(_1986_),
    .A2(_1989_),
    .B1(_1991_),
    .Y(_1992_));
 sky130_fd_sc_hs__a221oi_4 _7063_ (.A1(_1841_),
    .A2(_1976_),
    .B1(_1978_),
    .B2(_1874_),
    .C1(_1992_),
    .Y(_1993_));
 sky130_fd_sc_hs__nand2_1 _7064_ (.A(net198),
    .B(_1953_),
    .Y(_1994_));
 sky130_fd_sc_hs__a21oi_1 _7065_ (.A1(_1993_),
    .A2(_1994_),
    .B1(_1983_),
    .Y(_1995_));
 sky130_fd_sc_hs__a211o_2 _7066_ (.A1(_1328_),
    .A2(_0436_),
    .B1(_1380_),
    .C1(_1995_),
    .X(net332));
 sky130_fd_sc_hs__o21ai_1 _7067_ (.A1(_4040_),
    .A2(_1938_),
    .B1(_1773_),
    .Y(_1996_));
 sky130_fd_sc_hs__o2bb2ai_1 _7068_ (.A1_N(_4039_),
    .A2_N(_1938_),
    .B1(_1930_),
    .B2(_4041_),
    .Y(_1997_));
 sky130_fd_sc_hs__a21oi_2 _7069_ (.A1(_1768_),
    .A2(_1996_),
    .B1(_1997_),
    .Y(_1998_));
 sky130_fd_sc_hs__nor2_2 _7070_ (.A(_1734_),
    .B(_1967_),
    .Y(_1999_));
 sky130_fd_sc_hs__a211oi_4 _7071_ (.A1(_1890_),
    .A2(_1956_),
    .B1(_1860_),
    .C1(_1920_),
    .Y(_2000_));
 sky130_fd_sc_hs__a2111oi_4 _7072_ (.A1(net199),
    .A2(_1953_),
    .B1(_1998_),
    .C1(_1999_),
    .D1(_2000_),
    .Y(_2001_));
 sky130_fd_sc_hs__nand2_1 _7073_ (.A(_1606_),
    .B(_0446_),
    .Y(_2002_));
 sky130_fd_sc_hs__o211ai_4 _7074_ (.A1(_1937_),
    .A2(_2001_),
    .B1(_2002_),
    .C1(_1396_),
    .Y(net333));
 sky130_fd_sc_hs__o21ai_1 _7075_ (.A1(_4046_),
    .A2(_1938_),
    .B1(_1773_),
    .Y(_2003_));
 sky130_fd_sc_hs__o2bb2ai_1 _7076_ (.A1_N(_4045_),
    .A2_N(_1938_),
    .B1(_1930_),
    .B2(_4047_),
    .Y(_2004_));
 sky130_fd_sc_hs__a21oi_2 _7077_ (.A1(_1768_),
    .A2(_2003_),
    .B1(_2004_),
    .Y(_2005_));
 sky130_fd_sc_hs__o2bb2ai_4 _7078_ (.A1_N(_1874_),
    .A2_N(_1943_),
    .B1(_1949_),
    .B2(_1734_),
    .Y(_2006_));
 sky130_fd_sc_hs__a211oi_4 _7079_ (.A1(net200),
    .A2(_1840_),
    .B1(_2005_),
    .C1(_2006_),
    .Y(_2007_));
 sky130_fd_sc_hs__nand2_1 _7080_ (.A(_1606_),
    .B(_0449_),
    .Y(_2008_));
 sky130_fd_sc_hs__o211ai_4 _7081_ (.A1(_1937_),
    .A2(_2007_),
    .B1(_2008_),
    .C1(_1418_),
    .Y(net334));
 sky130_fd_sc_hs__buf_8 _7082_ (.A(_1241_),
    .X(_2009_));
 sky130_fd_sc_hs__nand2_1 _7083_ (.A(_4051_),
    .B(_1772_),
    .Y(_2010_));
 sky130_fd_sc_hs__o21ai_1 _7084_ (.A1(_4052_),
    .A2(_1771_),
    .B1(_1739_),
    .Y(_2011_));
 sky130_fd_sc_hs__nand2_1 _7085_ (.A(_1742_),
    .B(_2011_),
    .Y(_2012_));
 sky130_fd_sc_hs__o211ai_2 _7086_ (.A1(_4053_),
    .A2(_1930_),
    .B1(_2010_),
    .C1(_2012_),
    .Y(_2013_));
 sky130_fd_sc_hs__nand2_1 _7087_ (.A(_1835_),
    .B(_1919_),
    .Y(_2014_));
 sky130_fd_sc_hs__nand2_1 _7088_ (.A(net201),
    .B(_1928_),
    .Y(_2015_));
 sky130_fd_sc_hs__o2111a_1 _7089_ (.A1(_1734_),
    .A2(_1927_),
    .B1(_2013_),
    .C1(_2014_),
    .D1(_2015_),
    .X(_2016_));
 sky130_fd_sc_hs__nor2_1 _7090_ (.A(_1983_),
    .B(_2016_),
    .Y(_2017_));
 sky130_fd_sc_hs__a211o_2 _7091_ (.A1(_2009_),
    .A2(_0586_),
    .B1(_1425_),
    .C1(_2017_),
    .X(net335));
 sky130_fd_sc_hs__mux4_4 _7092_ (.A0(net41),
    .A1(net3),
    .A2(net24),
    .A3(net23),
    .S0(_1807_),
    .S1(_1808_),
    .X(_2018_));
 sky130_fd_sc_hs__mux2i_4 _7093_ (.A0(_1899_),
    .A1(_2018_),
    .S(_1758_),
    .Y(_2019_));
 sky130_fd_sc_hs__mux2i_4 _7094_ (.A0(_1945_),
    .A1(_2019_),
    .S(_1851_),
    .Y(_2020_));
 sky130_fd_sc_hs__mux4_4 _7095_ (.A0(net37),
    .A1(net38),
    .A2(net28),
    .A3(net27),
    .S0(_0596_),
    .S1(_1747_),
    .X(_2021_));
 sky130_fd_sc_hs__mux4_4 _7096_ (.A0(net39),
    .A1(net40),
    .A2(net26),
    .A3(net25),
    .S0(_1807_),
    .S1(_1808_),
    .X(_2022_));
 sky130_fd_sc_hs__mux2i_4 _7097_ (.A0(_2021_),
    .A1(_2022_),
    .S(_1794_),
    .Y(_2023_));
 sky130_fd_sc_hs__nand2_1 _7098_ (.A(_3933_),
    .B(_1819_),
    .Y(_2024_));
 sky130_fd_sc_hs__nand2_1 _7099_ (.A(_0596_),
    .B(_1816_),
    .Y(_2025_));
 sky130_fd_sc_hs__mux4_2 _7100_ (.A0(net35),
    .A1(net36),
    .A2(net30),
    .A3(net29),
    .S0(_1807_),
    .S1(_1808_),
    .X(_2026_));
 sky130_fd_sc_hs__and2_1 _7101_ (.A(_1794_),
    .B(_2026_),
    .X(_2027_));
 sky130_fd_sc_hs__a311oi_4 _7102_ (.A1(_1758_),
    .A2(_2024_),
    .A3(_2025_),
    .B1(_1806_),
    .C1(_2027_),
    .Y(_2028_));
 sky130_fd_sc_hs__a21oi_4 _7103_ (.A1(_1806_),
    .A2(_2023_),
    .B1(_2028_),
    .Y(_2029_));
 sky130_fd_sc_hs__mux2i_4 _7104_ (.A0(_2020_),
    .A1(_2029_),
    .S(_1844_),
    .Y(_2030_));
 sky130_fd_sc_hs__mux2i_4 _7105_ (.A0(_1956_),
    .A1(_2030_),
    .S(_1843_),
    .Y(_2031_));
 sky130_fd_sc_hs__a21oi_2 _7106_ (.A1(_1843_),
    .A2(_1961_),
    .B1(_1859_),
    .Y(_2032_));
 sky130_fd_sc_hs__o21ai_1 _7107_ (.A1(_3944_),
    .A2(_1775_),
    .B1(_1876_),
    .Y(_2033_));
 sky130_fd_sc_hs__o2bb2ai_1 _7108_ (.A1_N(_3943_),
    .A2_N(_1912_),
    .B1(_1777_),
    .B2(_3945_),
    .Y(_2034_));
 sky130_fd_sc_hs__a21oi_4 _7109_ (.A1(_1875_),
    .A2(_2033_),
    .B1(_2034_),
    .Y(_2035_));
 sky130_fd_sc_hs__a221o_1 _7110_ (.A1(net202),
    .A2(_1928_),
    .B1(_1748_),
    .B2(_2032_),
    .C1(_2035_),
    .X(_2036_));
 sky130_fd_sc_hs__a21oi_2 _7111_ (.A1(_1836_),
    .A2(_2031_),
    .B1(_2036_),
    .Y(_2037_));
 sky130_fd_sc_hs__a22o_2 _7112_ (.A1(_0447_),
    .A2(_1144_),
    .B1(_1719_),
    .B2(_3716_),
    .X(_2038_));
 sky130_fd_sc_hs__a22oi_4 _7113_ (.A1(_2009_),
    .A2(_0447_),
    .B1(_2038_),
    .B2(_0104_),
    .Y(_2039_));
 sky130_fd_sc_hs__o21ai_4 _7114_ (.A1(_1839_),
    .A2(_2037_),
    .B1(_2039_),
    .Y(net336));
 sky130_fd_sc_hs__o21ai_1 _7115_ (.A1(_4058_),
    .A2(_1775_),
    .B1(_1876_),
    .Y(_2040_));
 sky130_fd_sc_hs__o2bb2ai_1 _7116_ (.A1_N(_4057_),
    .A2_N(_1912_),
    .B1(_1777_),
    .B2(_4059_),
    .Y(_2041_));
 sky130_fd_sc_hs__a21oi_4 _7117_ (.A1(_1875_),
    .A2(_2040_),
    .B1(_2041_),
    .Y(_2042_));
 sky130_fd_sc_hs__a221o_1 _7118_ (.A1(_1874_),
    .A2(_1889_),
    .B1(_1910_),
    .B2(_1841_),
    .C1(_2042_),
    .X(_2043_));
 sky130_fd_sc_hs__a21oi_2 _7119_ (.A1(net203),
    .A2(_1840_),
    .B1(_2043_),
    .Y(_2044_));
 sky130_fd_sc_hs__a21oi_1 _7120_ (.A1(_1242_),
    .A2(_0588_),
    .B1(_1450_),
    .Y(_2045_));
 sky130_fd_sc_hs__o21ai_4 _7121_ (.A1(_1839_),
    .A2(_2044_),
    .B1(_2045_),
    .Y(net337));
 sky130_fd_sc_hs__o21ai_1 _7122_ (.A1(_4064_),
    .A2(_1912_),
    .B1(_1876_),
    .Y(_2046_));
 sky130_fd_sc_hs__o2bb2ai_1 _7123_ (.A1_N(_4063_),
    .A2_N(_1912_),
    .B1(_1777_),
    .B2(_4065_),
    .Y(_2047_));
 sky130_fd_sc_hs__a21oi_4 _7124_ (.A1(_1875_),
    .A2(_2046_),
    .B1(_2047_),
    .Y(_2048_));
 sky130_fd_sc_hs__a221oi_2 _7125_ (.A1(_1874_),
    .A2(_1861_),
    .B1(_1873_),
    .B2(_1841_),
    .C1(_2048_),
    .Y(_2049_));
 sky130_fd_sc_hs__nand2_1 _7126_ (.A(net204),
    .B(_1953_),
    .Y(_2050_));
 sky130_fd_sc_hs__a21oi_2 _7127_ (.A1(_2049_),
    .A2(_2050_),
    .B1(_1983_),
    .Y(_2051_));
 sky130_fd_sc_hs__a21oi_4 _7128_ (.A1(_1242_),
    .A2(net109),
    .B1(_2051_),
    .Y(_2052_));
 sky130_fd_sc_hs__nand2_8 _7129_ (.A(_1460_),
    .B(_2052_),
    .Y(net338));
 sky130_fd_sc_hs__o21ai_1 _7130_ (.A1(_4070_),
    .A2(_1938_),
    .B1(_1773_),
    .Y(_2053_));
 sky130_fd_sc_hs__o2bb2ai_1 _7131_ (.A1_N(_4069_),
    .A2_N(_1938_),
    .B1(_1930_),
    .B2(_4071_),
    .Y(_2054_));
 sky130_fd_sc_hs__a21oi_2 _7132_ (.A1(_1768_),
    .A2(_2053_),
    .B1(_2054_),
    .Y(_2055_));
 sky130_fd_sc_hs__a21oi_4 _7133_ (.A1(_1844_),
    .A2(_1954_),
    .B1(_1865_),
    .Y(_2056_));
 sky130_fd_sc_hs__nor2b_1 _7134_ (.A(_1803_),
    .B_N(_1955_),
    .Y(_2057_));
 sky130_fd_sc_hs__a211oi_4 _7135_ (.A1(_1862_),
    .A2(_2020_),
    .B1(_2057_),
    .C1(_1751_),
    .Y(_2058_));
 sky130_fd_sc_hs__a21oi_4 _7136_ (.A1(_1751_),
    .A2(_2056_),
    .B1(_2058_),
    .Y(_2059_));
 sky130_fd_sc_hs__nand2_2 _7137_ (.A(_1758_),
    .B(_1760_),
    .Y(_2060_));
 sky130_fd_sc_hs__mux2i_4 _7138_ (.A0(_1790_),
    .A1(_1765_),
    .S(_2060_),
    .Y(_2061_));
 sky130_fd_sc_hs__nor2_1 _7139_ (.A(_1805_),
    .B(_2061_),
    .Y(_2062_));
 sky130_fd_sc_hs__a21oi_4 _7140_ (.A1(_1862_),
    .A2(_1962_),
    .B1(_2062_),
    .Y(_2063_));
 sky130_fd_sc_hs__o21a_1 _7141_ (.A1(_1751_),
    .A2(_2063_),
    .B1(_1766_),
    .X(_2064_));
 sky130_fd_sc_hs__o2bb2ai_2 _7142_ (.A1_N(_1748_),
    .A2_N(_2059_),
    .B1(_2064_),
    .B2(_1920_),
    .Y(_2065_));
 sky130_fd_sc_hs__a211oi_4 _7143_ (.A1(net205),
    .A2(_1840_),
    .B1(_2055_),
    .C1(_2065_),
    .Y(_2066_));
 sky130_fd_sc_hs__a21oi_1 _7144_ (.A1(_1328_),
    .A2(_0520_),
    .B1(_1477_),
    .Y(_2067_));
 sky130_fd_sc_hs__o21ai_4 _7145_ (.A1(_1839_),
    .A2(_2066_),
    .B1(_2067_),
    .Y(net339));
 sky130_fd_sc_hs__a21oi_4 _7146_ (.A1(_1805_),
    .A2(_1795_),
    .B1(_1865_),
    .Y(_2068_));
 sky130_fd_sc_hs__nor2b_2 _7147_ (.A(_1756_),
    .B_N(_1802_),
    .Y(_2069_));
 sky130_fd_sc_hs__a211oi_4 _7148_ (.A1(_1844_),
    .A2(_1831_),
    .B1(_2069_),
    .C1(_1750_),
    .Y(_2070_));
 sky130_fd_sc_hs__a21oi_4 _7149_ (.A1(_1751_),
    .A2(_2068_),
    .B1(_2070_),
    .Y(_2071_));
 sky130_fd_sc_hs__o21ai_2 _7150_ (.A1(_0596_),
    .A2(_2060_),
    .B1(_1762_),
    .Y(_2072_));
 sky130_fd_sc_hs__nor2_1 _7151_ (.A(_1754_),
    .B(_1805_),
    .Y(_2073_));
 sky130_fd_sc_hs__a22oi_4 _7152_ (.A1(_1844_),
    .A2(_1973_),
    .B1(_2072_),
    .B2(_2073_),
    .Y(_2074_));
 sky130_fd_sc_hs__a21oi_4 _7153_ (.A1(_1843_),
    .A2(_2074_),
    .B1(_1860_),
    .Y(_2075_));
 sky130_fd_sc_hs__o21ai_1 _7154_ (.A1(_4076_),
    .A2(_1987_),
    .B1(_1988_),
    .Y(_2076_));
 sky130_fd_sc_hs__o2bb2ai_1 _7155_ (.A1_N(_4075_),
    .A2_N(_1987_),
    .B1(_1990_),
    .B2(_4077_),
    .Y(_2077_));
 sky130_fd_sc_hs__a21oi_4 _7156_ (.A1(_1986_),
    .A2(_2076_),
    .B1(_2077_),
    .Y(_2078_));
 sky130_fd_sc_hs__a221oi_4 _7157_ (.A1(_1841_),
    .A2(_2071_),
    .B1(_2075_),
    .B2(_1874_),
    .C1(_2078_),
    .Y(_2079_));
 sky130_fd_sc_hs__nand2_1 _7158_ (.A(net206),
    .B(_1953_),
    .Y(_2080_));
 sky130_fd_sc_hs__a21oi_1 _7159_ (.A1(_2079_),
    .A2(_2080_),
    .B1(_1983_),
    .Y(_2081_));
 sky130_fd_sc_hs__a211o_4 _7160_ (.A1(_2009_),
    .A2(_0526_),
    .B1(_1499_),
    .C1(_2081_),
    .X(net340));
 sky130_fd_sc_hs__a21oi_2 _7161_ (.A1(_1843_),
    .A2(_2068_),
    .B1(_1860_),
    .Y(_2082_));
 sky130_fd_sc_hs__nand2_1 _7162_ (.A(_1836_),
    .B(_2082_),
    .Y(_2083_));
 sky130_fd_sc_hs__nand2b_1 _7163_ (.A_N(_1862_),
    .B(_1974_),
    .Y(_2084_));
 sky130_fd_sc_hs__mux2i_4 _7164_ (.A0(_2018_),
    .A1(_2022_),
    .S(_1757_),
    .Y(_2085_));
 sky130_fd_sc_hs__nand2_1 _7165_ (.A(_1885_),
    .B(_2085_),
    .Y(_2086_));
 sky130_fd_sc_hs__o211ai_1 _7166_ (.A1(_1885_),
    .A2(_1901_),
    .B1(_2086_),
    .C1(_1862_),
    .Y(_2087_));
 sky130_fd_sc_hs__nand3_4 _7167_ (.A(_1890_),
    .B(_2084_),
    .C(_2087_),
    .Y(_2088_));
 sky130_fd_sc_hs__nand2_2 _7168_ (.A(_1751_),
    .B(_2074_),
    .Y(_2089_));
 sky130_fd_sc_hs__clkbuf_4 _7169_ (.A(_1771_),
    .X(_2090_));
 sky130_fd_sc_hs__o21ai_1 _7170_ (.A1(_4082_),
    .A2(_2090_),
    .B1(_1739_),
    .Y(_2091_));
 sky130_fd_sc_hs__o2bb2ai_1 _7171_ (.A1_N(_4081_),
    .A2_N(_1771_),
    .B1(_1776_),
    .B2(_4083_),
    .Y(_2092_));
 sky130_fd_sc_hs__a21oi_2 _7172_ (.A1(_1742_),
    .A2(_2091_),
    .B1(_2092_),
    .Y(_2093_));
 sky130_fd_sc_hs__a31oi_2 _7173_ (.A1(_1841_),
    .A2(_2088_),
    .A3(_2089_),
    .B1(_2093_),
    .Y(_2094_));
 sky130_fd_sc_hs__nand2_1 _7174_ (.A(net207),
    .B(_1953_),
    .Y(_2095_));
 sky130_fd_sc_hs__a31oi_4 _7175_ (.A1(_2083_),
    .A2(_2094_),
    .A3(_2095_),
    .B1(_1744_),
    .Y(_2096_));
 sky130_fd_sc_hs__a211o_2 _7176_ (.A1(_2009_),
    .A2(_0527_),
    .B1(_1518_),
    .C1(_2096_),
    .X(net341));
 sky130_fd_sc_hs__a21oi_4 _7177_ (.A1(_1843_),
    .A2(_2056_),
    .B1(_1860_),
    .Y(_2097_));
 sky130_fd_sc_hs__mux2i_4 _7178_ (.A0(_1810_),
    .A1(_1825_),
    .S(_1822_),
    .Y(_2098_));
 sky130_fd_sc_hs__mux2i_4 _7179_ (.A0(_1869_),
    .A1(_2098_),
    .S(_1885_),
    .Y(_2099_));
 sky130_fd_sc_hs__mux2i_4 _7180_ (.A0(_1965_),
    .A1(_2099_),
    .S(_1844_),
    .Y(_2100_));
 sky130_fd_sc_hs__mux2i_4 _7181_ (.A0(_2063_),
    .A1(_2100_),
    .S(_1843_),
    .Y(_2101_));
 sky130_fd_sc_hs__o21ai_1 _7182_ (.A1(_4088_),
    .A2(_1987_),
    .B1(_1988_),
    .Y(_2102_));
 sky130_fd_sc_hs__o2bb2ai_1 _7183_ (.A1_N(_4087_),
    .A2_N(_1987_),
    .B1(_1990_),
    .B2(_4089_),
    .Y(_2103_));
 sky130_fd_sc_hs__a21oi_4 _7184_ (.A1(_1986_),
    .A2(_2102_),
    .B1(_2103_),
    .Y(_2104_));
 sky130_fd_sc_hs__a221oi_4 _7185_ (.A1(_1835_),
    .A2(_2097_),
    .B1(_2101_),
    .B2(_1841_),
    .C1(_2104_),
    .Y(_2105_));
 sky130_fd_sc_hs__nand2_1 _7186_ (.A(net208),
    .B(_1953_),
    .Y(_2106_));
 sky130_fd_sc_hs__a21oi_1 _7187_ (.A1(_2105_),
    .A2(_2106_),
    .B1(_1983_),
    .Y(_2107_));
 sky130_fd_sc_hs__a211o_2 _7188_ (.A1(_2009_),
    .A2(_0529_),
    .B1(_1539_),
    .C1(_2107_),
    .X(net342));
 sky130_fd_sc_hs__mux2i_4 _7189_ (.A0(_2019_),
    .A1(_2023_),
    .S(_1851_),
    .Y(_2108_));
 sky130_fd_sc_hs__mux2i_4 _7190_ (.A0(_1947_),
    .A1(_2108_),
    .S(_1805_),
    .Y(_2109_));
 sky130_fd_sc_hs__mux2i_4 _7191_ (.A0(_1858_),
    .A1(_2109_),
    .S(_1842_),
    .Y(_2110_));
 sky130_fd_sc_hs__a21oi_4 _7192_ (.A1(_1890_),
    .A2(_1866_),
    .B1(_1860_),
    .Y(_2111_));
 sky130_fd_sc_hs__o21ai_1 _7193_ (.A1(_4094_),
    .A2(_2090_),
    .B1(_1988_),
    .Y(_2112_));
 sky130_fd_sc_hs__o2bb2ai_1 _7194_ (.A1_N(_4093_),
    .A2_N(_2090_),
    .B1(_1990_),
    .B2(_4095_),
    .Y(_2113_));
 sky130_fd_sc_hs__a21oi_1 _7195_ (.A1(_1986_),
    .A2(_2112_),
    .B1(_2113_),
    .Y(_2114_));
 sky130_fd_sc_hs__a221o_2 _7196_ (.A1(_1747_),
    .A2(_2110_),
    .B1(_2111_),
    .B2(_1835_),
    .C1(_2114_),
    .X(_2115_));
 sky130_fd_sc_hs__a21oi_4 _7197_ (.A1(net209),
    .A2(_1840_),
    .B1(_2115_),
    .Y(_2116_));
 sky130_fd_sc_hs__nand2_1 _7198_ (.A(_1606_),
    .B(_0565_),
    .Y(_2117_));
 sky130_fd_sc_hs__o211ai_4 _7199_ (.A1(_1937_),
    .A2(_2116_),
    .B1(_2117_),
    .C1(_1557_),
    .Y(net343));
 sky130_fd_sc_hs__nand2_1 _7200_ (.A(_1885_),
    .B(_1811_),
    .Y(_2118_));
 sky130_fd_sc_hs__nand2_1 _7201_ (.A(_1806_),
    .B(_1827_),
    .Y(_2119_));
 sky130_fd_sc_hs__nor2b_1 _7202_ (.A(_1805_),
    .B_N(_1923_),
    .Y(_2120_));
 sky130_fd_sc_hs__a311oi_4 _7203_ (.A1(_1862_),
    .A2(_2118_),
    .A3(_2119_),
    .B1(_2120_),
    .C1(_1751_),
    .Y(_2121_));
 sky130_fd_sc_hs__a21oi_4 _7204_ (.A1(_1751_),
    .A2(_1888_),
    .B1(_2121_),
    .Y(_2122_));
 sky130_fd_sc_hs__and2_2 _7205_ (.A(_1842_),
    .B(_1803_),
    .X(_2123_));
 sky130_fd_sc_hs__mux2i_4 _7206_ (.A0(_1765_),
    .A1(_1908_),
    .S(_2123_),
    .Y(_2124_));
 sky130_fd_sc_hs__o21ai_1 _7207_ (.A1(_4100_),
    .A2(_1912_),
    .B1(_1876_),
    .Y(_2125_));
 sky130_fd_sc_hs__o2bb2ai_1 _7208_ (.A1_N(_4099_),
    .A2_N(_1987_),
    .B1(_1990_),
    .B2(_4101_),
    .Y(_2126_));
 sky130_fd_sc_hs__a21oi_4 _7209_ (.A1(_1875_),
    .A2(_2125_),
    .B1(_2126_),
    .Y(_2127_));
 sky130_fd_sc_hs__o21bai_1 _7210_ (.A1(_1920_),
    .A2(_2124_),
    .B1_N(_2127_),
    .Y(_2128_));
 sky130_fd_sc_hs__a221oi_4 _7211_ (.A1(net210),
    .A2(_1953_),
    .B1(_1748_),
    .B2(_2122_),
    .C1(_2128_),
    .Y(_2129_));
 sky130_fd_sc_hs__nand2_1 _7212_ (.A(_1606_),
    .B(_0566_),
    .Y(_2130_));
 sky130_fd_sc_hs__o211ai_4 _7213_ (.A1(_1937_),
    .A2(_2129_),
    .B1(_2130_),
    .C1(_1575_),
    .Y(net344));
 sky130_fd_sc_hs__mux2_1 _7214_ (.A0(_2026_),
    .A1(_2021_),
    .S(_1822_),
    .X(_2131_));
 sky130_fd_sc_hs__nand2_1 _7215_ (.A(_1806_),
    .B(_2085_),
    .Y(_2132_));
 sky130_fd_sc_hs__o211ai_1 _7216_ (.A1(_1806_),
    .A2(_2131_),
    .B1(_2132_),
    .C1(_1803_),
    .Y(_2133_));
 sky130_fd_sc_hs__o211ai_2 _7217_ (.A1(_1805_),
    .A2(_1903_),
    .B1(_2133_),
    .C1(_1842_),
    .Y(_2134_));
 sky130_fd_sc_hs__a21boi_4 _7218_ (.A1(_1750_),
    .A2(_1918_),
    .B1_N(_2134_),
    .Y(_2135_));
 sky130_fd_sc_hs__a21oi_2 _7219_ (.A1(_1885_),
    .A2(_2123_),
    .B1(_1765_),
    .Y(_2136_));
 sky130_fd_sc_hs__a31oi_4 _7220_ (.A1(_1885_),
    .A2(_1886_),
    .A3(_2123_),
    .B1(_2136_),
    .Y(_2137_));
 sky130_fd_sc_hs__o21ai_1 _7221_ (.A1(_4106_),
    .A2(_2090_),
    .B1(_1988_),
    .Y(_2138_));
 sky130_fd_sc_hs__o2bb2ai_1 _7222_ (.A1_N(_4105_),
    .A2_N(_2090_),
    .B1(_1990_),
    .B2(_4107_),
    .Y(_2139_));
 sky130_fd_sc_hs__a21oi_1 _7223_ (.A1(_1986_),
    .A2(_2138_),
    .B1(_2139_),
    .Y(_2140_));
 sky130_fd_sc_hs__a221o_2 _7224_ (.A1(_1747_),
    .A2(_2135_),
    .B1(_2137_),
    .B2(_1835_),
    .C1(_2140_),
    .X(_2141_));
 sky130_fd_sc_hs__a21oi_2 _7225_ (.A1(net211),
    .A2(_1840_),
    .B1(_2141_),
    .Y(_2142_));
 sky130_fd_sc_hs__nand2_1 _7226_ (.A(_1606_),
    .B(net111),
    .Y(_2143_));
 sky130_fd_sc_hs__o211ai_4 _7227_ (.A1(_1937_),
    .A2(_2142_),
    .B1(_2143_),
    .C1(_1598_),
    .Y(net345));
 sky130_fd_sc_hs__and2_1 _7228_ (.A(_1822_),
    .B(_1809_),
    .X(_2144_));
 sky130_fd_sc_hs__a211oi_4 _7229_ (.A1(_1758_),
    .A2(_1817_),
    .B1(_2144_),
    .C1(_1787_),
    .Y(_2145_));
 sky130_fd_sc_hs__a21oi_4 _7230_ (.A1(_1806_),
    .A2(_2098_),
    .B1(_2145_),
    .Y(_2146_));
 sky130_fd_sc_hs__nor2b_1 _7231_ (.A(_1756_),
    .B_N(_1871_),
    .Y(_2147_));
 sky130_fd_sc_hs__a211oi_4 _7232_ (.A1(_1844_),
    .A2(_2146_),
    .B1(_2147_),
    .C1(_1750_),
    .Y(_2148_));
 sky130_fd_sc_hs__a21oi_4 _7233_ (.A1(_1751_),
    .A2(_1942_),
    .B1(_2148_),
    .Y(_2149_));
 sky130_fd_sc_hs__nand2_2 _7234_ (.A(_1890_),
    .B(_1944_),
    .Y(_2150_));
 sky130_fd_sc_hs__nand2_4 _7235_ (.A(_1766_),
    .B(_2150_),
    .Y(_2151_));
 sky130_fd_sc_hs__o21ai_1 _7236_ (.A1(_4112_),
    .A2(_1987_),
    .B1(_1988_),
    .Y(_2152_));
 sky130_fd_sc_hs__o2bb2ai_1 _7237_ (.A1_N(_4111_),
    .A2_N(_2090_),
    .B1(_1990_),
    .B2(_4113_),
    .Y(_2153_));
 sky130_fd_sc_hs__a21oi_4 _7238_ (.A1(_1986_),
    .A2(_2152_),
    .B1(_2153_),
    .Y(_2154_));
 sky130_fd_sc_hs__a221oi_4 _7239_ (.A1(_1747_),
    .A2(_2149_),
    .B1(_2151_),
    .B2(_1874_),
    .C1(_2154_),
    .Y(_2155_));
 sky130_fd_sc_hs__nand2_1 _7240_ (.A(net10),
    .B(_1953_),
    .Y(_2156_));
 sky130_fd_sc_hs__a21oi_1 _7241_ (.A1(_2155_),
    .A2(_2156_),
    .B1(_1983_),
    .Y(_2157_));
 sky130_fd_sc_hs__a211o_2 _7242_ (.A1(_2009_),
    .A2(net112),
    .B1(_1627_),
    .C1(_2157_),
    .X(net346));
 sky130_fd_sc_hs__o21ai_1 _7243_ (.A1(_3950_),
    .A2(_1775_),
    .B1(_1876_),
    .Y(_2158_));
 sky130_fd_sc_hs__o2bb2ai_1 _7244_ (.A1_N(_3949_),
    .A2_N(_1912_),
    .B1(_1777_),
    .B2(_3951_),
    .Y(_2159_));
 sky130_fd_sc_hs__a21oi_4 _7245_ (.A1(_1875_),
    .A2(_2158_),
    .B1(_2159_),
    .Y(_2160_));
 sky130_fd_sc_hs__a221o_1 _7246_ (.A1(net213),
    .A2(_1928_),
    .B1(_1748_),
    .B2(_2151_),
    .C1(_2160_),
    .X(_2161_));
 sky130_fd_sc_hs__a21oi_2 _7247_ (.A1(_1836_),
    .A2(_2149_),
    .B1(_2161_),
    .Y(_2162_));
 sky130_fd_sc_hs__nand2_1 _7248_ (.A(_3718_),
    .B(_1719_),
    .Y(_2163_));
 sky130_fd_sc_hs__nand2_2 _7249_ (.A(_1145_),
    .B(_2163_),
    .Y(_2164_));
 sky130_fd_sc_hs__a22oi_4 _7250_ (.A1(_2009_),
    .A2(_0450_),
    .B1(_2164_),
    .B2(_0104_),
    .Y(_2165_));
 sky130_fd_sc_hs__o21ai_4 _7251_ (.A1(_1839_),
    .A2(_2162_),
    .B1(_2165_),
    .Y(net347));
 sky130_fd_sc_hs__o21ai_1 _7252_ (.A1(_4118_),
    .A2(_2090_),
    .B1(_1988_),
    .Y(_2166_));
 sky130_fd_sc_hs__o2bb2ai_1 _7253_ (.A1_N(_4117_),
    .A2_N(_1771_),
    .B1(_1990_),
    .B2(_4119_),
    .Y(_2167_));
 sky130_fd_sc_hs__a21oi_2 _7254_ (.A1(_1986_),
    .A2(_2166_),
    .B1(_2167_),
    .Y(_2168_));
 sky130_fd_sc_hs__a221o_2 _7255_ (.A1(_1835_),
    .A2(_2032_),
    .B1(_2031_),
    .B2(_1747_),
    .C1(_2168_),
    .X(_2169_));
 sky130_fd_sc_hs__a21oi_2 _7256_ (.A1(net214),
    .A2(_1840_),
    .B1(_2169_),
    .Y(_2170_));
 sky130_fd_sc_hs__nand2_1 _7257_ (.A(_1606_),
    .B(_0567_),
    .Y(_2171_));
 sky130_fd_sc_hs__o211ai_4 _7258_ (.A1(_1983_),
    .A2(_2170_),
    .B1(_2171_),
    .C1(_1638_),
    .Y(net348));
 sky130_fd_sc_hs__o21ai_1 _7259_ (.A1(_3930_),
    .A2(_1987_),
    .B1(_1988_),
    .Y(_2172_));
 sky130_fd_sc_hs__o2bb2ai_1 _7260_ (.A1_N(_3929_),
    .A2_N(_2090_),
    .B1(_1990_),
    .B2(_3931_),
    .Y(_2173_));
 sky130_fd_sc_hs__a21oi_2 _7261_ (.A1(_1986_),
    .A2(_2172_),
    .B1(_2173_),
    .Y(_2174_));
 sky130_fd_sc_hs__a221oi_4 _7262_ (.A1(_1747_),
    .A2(_1834_),
    .B1(_1874_),
    .B2(_1767_),
    .C1(_2174_),
    .Y(_2175_));
 sky130_fd_sc_hs__nand2_1 _7263_ (.A(net215),
    .B(_1953_),
    .Y(_2176_));
 sky130_fd_sc_hs__a21oi_2 _7264_ (.A1(_2175_),
    .A2(_2176_),
    .B1(_1983_),
    .Y(_2177_));
 sky130_fd_sc_hs__a211o_2 _7265_ (.A1(_2009_),
    .A2(_0382_),
    .B1(_1651_),
    .C1(_2177_),
    .X(net349));
 sky130_fd_sc_hs__o21ai_1 _7266_ (.A1(_3956_),
    .A2(_1775_),
    .B1(_1876_),
    .Y(_2178_));
 sky130_fd_sc_hs__o2bb2ai_1 _7267_ (.A1_N(_3955_),
    .A2_N(_1912_),
    .B1(_1777_),
    .B2(_3957_),
    .Y(_2179_));
 sky130_fd_sc_hs__a21oi_4 _7268_ (.A1(_1875_),
    .A2(_2178_),
    .B1(_2179_),
    .Y(_2180_));
 sky130_fd_sc_hs__a221o_1 _7269_ (.A1(net216),
    .A2(_1928_),
    .B1(_1748_),
    .B2(_2137_),
    .C1(_2180_),
    .X(_2181_));
 sky130_fd_sc_hs__a21oi_4 _7270_ (.A1(_1836_),
    .A2(_2135_),
    .B1(_2181_),
    .Y(_2182_));
 sky130_fd_sc_hs__a21oi_4 _7271_ (.A1(_1328_),
    .A2(_0572_),
    .B1(_1161_),
    .Y(_2183_));
 sky130_fd_sc_hs__o21ai_4 _7272_ (.A1(_1839_),
    .A2(_2182_),
    .B1(_2183_),
    .Y(net350));
 sky130_fd_sc_hs__o21ai_1 _7273_ (.A1(_3962_),
    .A2(_1772_),
    .B1(_1773_),
    .Y(_2184_));
 sky130_fd_sc_hs__o2bb2ai_1 _7274_ (.A1_N(_3961_),
    .A2_N(_1772_),
    .B1(_1930_),
    .B2(_3963_),
    .Y(_2185_));
 sky130_fd_sc_hs__a21oi_1 _7275_ (.A1(_1768_),
    .A2(_2184_),
    .B1(_2185_),
    .Y(_2186_));
 sky130_fd_sc_hs__a21oi_1 _7276_ (.A1(net217),
    .A2(_1928_),
    .B1(_2186_),
    .Y(_2187_));
 sky130_fd_sc_hs__o21ai_1 _7277_ (.A1(_1734_),
    .A2(_2124_),
    .B1(_2187_),
    .Y(_2188_));
 sky130_fd_sc_hs__a21oi_2 _7278_ (.A1(_1836_),
    .A2(_2122_),
    .B1(_2188_),
    .Y(_2189_));
 sky130_fd_sc_hs__nand2_1 _7279_ (.A(_3730_),
    .B(_1719_),
    .Y(_2190_));
 sky130_fd_sc_hs__nand2_4 _7280_ (.A(_1179_),
    .B(_2190_),
    .Y(_2191_));
 sky130_fd_sc_hs__a22oi_4 _7281_ (.A1(_2009_),
    .A2(_0573_),
    .B1(_2191_),
    .B2(_0104_),
    .Y(_2192_));
 sky130_fd_sc_hs__o21ai_4 _7282_ (.A1(_1839_),
    .A2(_2189_),
    .B1(_2192_),
    .Y(net351));
 sky130_fd_sc_hs__o21ai_1 _7283_ (.A1(_3968_),
    .A2(_1775_),
    .B1(_1876_),
    .Y(_2193_));
 sky130_fd_sc_hs__o2bb2ai_1 _7284_ (.A1_N(_3967_),
    .A2_N(_1912_),
    .B1(_1777_),
    .B2(_3969_),
    .Y(_2194_));
 sky130_fd_sc_hs__a21oi_2 _7285_ (.A1(_1875_),
    .A2(_2193_),
    .B1(_2194_),
    .Y(_2195_));
 sky130_fd_sc_hs__a221o_1 _7286_ (.A1(net218),
    .A2(_1928_),
    .B1(_1841_),
    .B2(_2111_),
    .C1(_2195_),
    .X(_2196_));
 sky130_fd_sc_hs__a21oi_2 _7287_ (.A1(_1836_),
    .A2(_2110_),
    .B1(_2196_),
    .Y(_2197_));
 sky130_fd_sc_hs__nand2_1 _7288_ (.A(_3739_),
    .B(_1719_),
    .Y(_2198_));
 sky130_fd_sc_hs__nand2_4 _7289_ (.A(_1187_),
    .B(_2198_),
    .Y(_2199_));
 sky130_fd_sc_hs__a22oi_4 _7290_ (.A1(_2009_),
    .A2(_0574_),
    .B1(_2199_),
    .B2(_0104_),
    .Y(_2200_));
 sky130_fd_sc_hs__o21ai_4 _7291_ (.A1(_1937_),
    .A2(_2197_),
    .B1(_2200_),
    .Y(net352));
 sky130_fd_sc_hs__o21ai_1 _7292_ (.A1(_3974_),
    .A2(_1775_),
    .B1(_1876_),
    .Y(_2201_));
 sky130_fd_sc_hs__o2bb2ai_1 _7293_ (.A1_N(_3973_),
    .A2_N(_1912_),
    .B1(_1777_),
    .B2(_3975_),
    .Y(_2202_));
 sky130_fd_sc_hs__a21oi_4 _7294_ (.A1(_1875_),
    .A2(_2201_),
    .B1(_2202_),
    .Y(_2203_));
 sky130_fd_sc_hs__a221o_1 _7295_ (.A1(net219),
    .A2(_1928_),
    .B1(_1874_),
    .B2(_2101_),
    .C1(_2203_),
    .X(_2204_));
 sky130_fd_sc_hs__a21oi_2 _7296_ (.A1(_1748_),
    .A2(_2097_),
    .B1(_2204_),
    .Y(_2205_));
 sky130_fd_sc_hs__a21oi_1 _7297_ (.A1(_1328_),
    .A2(_0575_),
    .B1(_1204_),
    .Y(_2206_));
 sky130_fd_sc_hs__o21ai_4 _7298_ (.A1(_1937_),
    .A2(_2205_),
    .B1(_2206_),
    .Y(net353));
 sky130_fd_sc_hs__o21ai_1 _7299_ (.A1(_3980_),
    .A2(_1987_),
    .B1(_1988_),
    .Y(_2207_));
 sky130_fd_sc_hs__o2bb2ai_1 _7300_ (.A1_N(_3979_),
    .A2_N(_2090_),
    .B1(_1990_),
    .B2(_3981_),
    .Y(_2208_));
 sky130_fd_sc_hs__a21oi_4 _7301_ (.A1(_1986_),
    .A2(_2207_),
    .B1(_2208_),
    .Y(_2209_));
 sky130_fd_sc_hs__a221o_1 _7302_ (.A1(net220),
    .A2(_1737_),
    .B1(_1841_),
    .B2(_2082_),
    .C1(_2209_),
    .X(_2210_));
 sky130_fd_sc_hs__a31oi_4 _7303_ (.A1(_1836_),
    .A2(_2088_),
    .A3(_2089_),
    .B1(_2210_),
    .Y(_2211_));
 sky130_fd_sc_hs__a21oi_2 _7304_ (.A1(_1328_),
    .A2(_0576_),
    .B1(_1217_),
    .Y(_2212_));
 sky130_fd_sc_hs__o21ai_4 _7305_ (.A1(_1937_),
    .A2(_2211_),
    .B1(_2212_),
    .Y(net354));
 sky130_fd_sc_hs__o21ai_1 _7306_ (.A1(_3986_),
    .A2(_2090_),
    .B1(_1988_),
    .Y(_2213_));
 sky130_fd_sc_hs__o2bb2ai_1 _7307_ (.A1_N(_3985_),
    .A2_N(_1771_),
    .B1(_1776_),
    .B2(_3987_),
    .Y(_2214_));
 sky130_fd_sc_hs__a21oi_2 _7308_ (.A1(_1986_),
    .A2(_2213_),
    .B1(_2214_),
    .Y(_2215_));
 sky130_fd_sc_hs__a221o_2 _7309_ (.A1(_1835_),
    .A2(_2071_),
    .B1(_2075_),
    .B2(_1747_),
    .C1(_2215_),
    .X(_2216_));
 sky130_fd_sc_hs__a21oi_2 _7310_ (.A1(net221),
    .A2(_1840_),
    .B1(_2216_),
    .Y(_2217_));
 sky130_fd_sc_hs__nand2_1 _7311_ (.A(_1606_),
    .B(_0577_),
    .Y(_2218_));
 sky130_fd_sc_hs__o211ai_4 _7312_ (.A1(_1983_),
    .A2(_2217_),
    .B1(_2218_),
    .C1(_1234_),
    .Y(net355));
 sky130_fd_sc_hs__o21ai_1 _7313_ (.A1(_3992_),
    .A2(_1772_),
    .B1(_1773_),
    .Y(_2219_));
 sky130_fd_sc_hs__o2bb2ai_1 _7314_ (.A1_N(_3991_),
    .A2_N(_1772_),
    .B1(_1930_),
    .B2(_3993_),
    .Y(_2220_));
 sky130_fd_sc_hs__a21oi_2 _7315_ (.A1(_1768_),
    .A2(_2219_),
    .B1(_2220_),
    .Y(_2221_));
 sky130_fd_sc_hs__a21oi_2 _7316_ (.A1(net222),
    .A2(_1928_),
    .B1(_2221_),
    .Y(_2222_));
 sky130_fd_sc_hs__o21ai_1 _7317_ (.A1(_1734_),
    .A2(_2064_),
    .B1(_2222_),
    .Y(_2223_));
 sky130_fd_sc_hs__a21oi_2 _7318_ (.A1(_1836_),
    .A2(_2059_),
    .B1(_2223_),
    .Y(_2224_));
 sky130_fd_sc_hs__a21oi_4 _7319_ (.A1(_1328_),
    .A2(_0578_),
    .B1(_1255_),
    .Y(_2225_));
 sky130_fd_sc_hs__o21ai_4 _7320_ (.A1(_1937_),
    .A2(_2224_),
    .B1(_2225_),
    .Y(net356));
 sky130_fd_sc_hs__fa_4 _7321_ (.A(_2226_),
    .B(_2227_),
    .CIN(_2228_),
    .COUT(_2229_),
    .SUM(net191));
 sky130_fd_sc_hs__fa_1 _7322_ (.A(_2230_),
    .B(_2231_),
    .CIN(_2232_),
    .COUT(_2233_),
    .SUM(_2234_));
 sky130_fd_sc_hs__fa_1 _7323_ (.A(_2235_),
    .B(_2236_),
    .CIN(_2237_),
    .COUT(_2238_),
    .SUM(_2239_));
 sky130_fd_sc_hs__fa_1 _7324_ (.A(_2240_),
    .B(_2241_),
    .CIN(_2242_),
    .COUT(_2243_),
    .SUM(_2244_));
 sky130_fd_sc_hs__fa_1 _7325_ (.A(_2245_),
    .B(_2246_),
    .CIN(_2247_),
    .COUT(_2248_),
    .SUM(_2249_));
 sky130_fd_sc_hs__fa_1 _7326_ (.A(_2250_),
    .B(_2238_),
    .CIN(_2251_),
    .COUT(_2252_),
    .SUM(_2253_));
 sky130_fd_sc_hs__fa_1 _7327_ (.A(_2254_),
    .B(_2255_),
    .CIN(_2256_),
    .COUT(_2257_),
    .SUM(_2258_));
 sky130_fd_sc_hs__fa_1 _7328_ (.A(_2259_),
    .B(_2260_),
    .CIN(_2261_),
    .COUT(_2262_),
    .SUM(_2263_));
 sky130_fd_sc_hs__fa_1 _7329_ (.A(_2264_),
    .B(_2265_),
    .CIN(_2266_),
    .COUT(_2267_),
    .SUM(_2268_));
 sky130_fd_sc_hs__fa_1 _7330_ (.A(_2269_),
    .B(_2270_),
    .CIN(_2271_),
    .COUT(_2272_),
    .SUM(_2273_));
 sky130_fd_sc_hs__fa_1 _7331_ (.A(_2274_),
    .B(_2275_),
    .CIN(_2276_),
    .COUT(_2277_),
    .SUM(_2278_));
 sky130_fd_sc_hs__fa_2 _7332_ (.A(_2279_),
    .B(_2280_),
    .CIN(_2281_),
    .COUT(_2282_),
    .SUM(_2283_));
 sky130_fd_sc_hs__fa_1 _7333_ (.A(_2283_),
    .B(_2284_),
    .CIN(_2285_),
    .COUT(_2286_),
    .SUM(_2287_));
 sky130_fd_sc_hs__fa_1 _7334_ (.A(_2288_),
    .B(_2267_),
    .CIN(_2287_),
    .COUT(_2289_),
    .SUM(_2290_));
 sky130_fd_sc_hs__fa_1 _7335_ (.A(_2291_),
    .B(_2292_),
    .CIN(_2293_),
    .COUT(_2294_),
    .SUM(_2295_));
 sky130_fd_sc_hs__fa_1 _7336_ (.A(_2296_),
    .B(_2297_),
    .CIN(_2298_),
    .COUT(_2299_),
    .SUM(_2300_));
 sky130_fd_sc_hs__fa_1 _7337_ (.A(_2301_),
    .B(_2302_),
    .CIN(_2303_),
    .COUT(_2304_),
    .SUM(_2305_));
 sky130_fd_sc_hs__fa_1 _7338_ (.A(_2306_),
    .B(_2286_),
    .CIN(_2305_),
    .COUT(_2307_),
    .SUM(_2308_));
 sky130_fd_sc_hs__fa_1 _7339_ (.A(_2309_),
    .B(_2289_),
    .CIN(_2308_),
    .COUT(_2310_),
    .SUM(_2311_));
 sky130_fd_sc_hs__fa_1 _7340_ (.A(_2313_),
    .B(_2314_),
    .CIN(_2315_),
    .COUT(_2316_),
    .SUM(_2317_));
 sky130_fd_sc_hs__fa_1 _7341_ (.A(_2318_),
    .B(_2319_),
    .CIN(_2320_),
    .COUT(_2321_),
    .SUM(_2322_));
 sky130_fd_sc_hs__fa_1 _7342_ (.A(_2323_),
    .B(_2324_),
    .CIN(_2325_),
    .COUT(_2326_),
    .SUM(_2327_));
 sky130_fd_sc_hs__fa_1 _7343_ (.A(_2328_),
    .B(_2329_),
    .CIN(_2330_),
    .COUT(_2331_),
    .SUM(_2332_));
 sky130_fd_sc_hs__fa_1 _7344_ (.A(_2333_),
    .B(_2332_),
    .CIN(_2299_),
    .COUT(_2334_),
    .SUM(_2335_));
 sky130_fd_sc_hs__fa_1 _7345_ (.A(_2336_),
    .B(_2304_),
    .CIN(_2327_),
    .COUT(_2337_),
    .SUM(_2338_));
 sky130_fd_sc_hs__fa_1 _7346_ (.A(_2339_),
    .B(_2307_),
    .CIN(_2338_),
    .COUT(_2340_),
    .SUM(_2341_));
 sky130_fd_sc_hs__fa_2 _7347_ (.A(_2343_),
    .B(_2344_),
    .CIN(_2345_),
    .COUT(_2346_),
    .SUM(_2347_));
 sky130_fd_sc_hs__fa_1 _7348_ (.A(_2348_),
    .B(_2349_),
    .CIN(_2350_),
    .COUT(_2351_),
    .SUM(_2352_));
 sky130_fd_sc_hs__fa_1 _7349_ (.A(_2353_),
    .B(_2354_),
    .CIN(_2355_),
    .COUT(_2356_),
    .SUM(_2357_));
 sky130_fd_sc_hs__fa_2 _7350_ (.A(_2358_),
    .B(_2359_),
    .CIN(_2360_),
    .COUT(_2361_),
    .SUM(_2362_));
 sky130_fd_sc_hs__fa_1 _7351_ (.A(_2363_),
    .B(_2364_),
    .CIN(_2365_),
    .COUT(_2366_),
    .SUM(_2367_));
 sky130_fd_sc_hs__fa_1 _7352_ (.A(_2331_),
    .B(_2367_),
    .CIN(_2321_),
    .COUT(_2368_),
    .SUM(_2369_));
 sky130_fd_sc_hs__fa_1 _7353_ (.A(_2370_),
    .B(_2326_),
    .CIN(_2362_),
    .COUT(_2371_),
    .SUM(_2372_));
 sky130_fd_sc_hs__fa_1 _7354_ (.A(_2373_),
    .B(_2337_),
    .CIN(_2372_),
    .COUT(_2374_),
    .SUM(_2375_));
 sky130_fd_sc_hs__fa_1 _7355_ (.A(_2376_),
    .B(_2377_),
    .CIN(_2378_),
    .COUT(_2379_),
    .SUM(_2380_));
 sky130_fd_sc_hs__fa_1 _7356_ (.A(_2381_),
    .B(_2382_),
    .CIN(_2383_),
    .COUT(_2384_),
    .SUM(_2385_));
 sky130_fd_sc_hs__fa_1 _7357_ (.A(_2386_),
    .B(_2387_),
    .CIN(_2388_),
    .COUT(_2389_),
    .SUM(_2390_));
 sky130_fd_sc_hs__fa_1 _7358_ (.A(_2391_),
    .B(_2392_),
    .CIN(_2393_),
    .COUT(_2394_),
    .SUM(_2395_));
 sky130_fd_sc_hs__fa_1 _7359_ (.A(_2366_),
    .B(_2395_),
    .CIN(_2356_),
    .COUT(_2396_),
    .SUM(_2397_));
 sky130_fd_sc_hs__fa_1 _7360_ (.A(_2398_),
    .B(_2361_),
    .CIN(_2390_),
    .COUT(_2399_),
    .SUM(_2400_));
 sky130_fd_sc_hs__fa_1 _7361_ (.A(_2401_),
    .B(_2371_),
    .CIN(_2400_),
    .COUT(_2402_),
    .SUM(_2403_));
 sky130_fd_sc_hs__fa_1 _7362_ (.A(_2404_),
    .B(_2374_),
    .CIN(_2403_),
    .COUT(_2405_),
    .SUM(_2406_));
 sky130_fd_sc_hs__fa_1 _7363_ (.A(_2408_),
    .B(_2409_),
    .CIN(_2410_),
    .COUT(_2411_),
    .SUM(_2412_));
 sky130_fd_sc_hs__fa_1 _7364_ (.A(_2413_),
    .B(_2414_),
    .CIN(_2415_),
    .COUT(_2416_),
    .SUM(_2417_));
 sky130_fd_sc_hs__fa_1 _7365_ (.A(_2418_),
    .B(_2419_),
    .CIN(_2420_),
    .COUT(_2421_),
    .SUM(_2422_));
 sky130_fd_sc_hs__fa_1 _7366_ (.A(_2423_),
    .B(_2424_),
    .CIN(_2425_),
    .COUT(_2426_),
    .SUM(_2427_));
 sky130_fd_sc_hs__fa_1 _7367_ (.A(_2428_),
    .B(_2429_),
    .CIN(_2430_),
    .COUT(_2431_),
    .SUM(_2432_));
 sky130_fd_sc_hs__fa_1 _7368_ (.A(_2432_),
    .B(_2389_),
    .CIN(_2422_),
    .COUT(_2433_),
    .SUM(_2434_));
 sky130_fd_sc_hs__fa_1 _7369_ (.A(_2435_),
    .B(_2436_),
    .CIN(_2437_),
    .COUT(_2438_),
    .SUM(_2439_));
 sky130_fd_sc_hs__fa_1 _7370_ (.A(_2440_),
    .B(_2399_),
    .CIN(_2434_),
    .COUT(_2441_),
    .SUM(_2442_));
 sky130_fd_sc_hs__fa_1 _7371_ (.A(_2443_),
    .B(_2402_),
    .CIN(_2442_),
    .COUT(_2444_),
    .SUM(_2445_));
 sky130_fd_sc_hs__fa_1 _7372_ (.A(_2446_),
    .B(_2447_),
    .CIN(_2448_),
    .COUT(_2449_),
    .SUM(_2450_));
 sky130_fd_sc_hs__fa_1 _7373_ (.A(_2451_),
    .B(_2452_),
    .CIN(_2453_),
    .COUT(_2454_),
    .SUM(_2455_));
 sky130_fd_sc_hs__fa_1 _7374_ (.A(_2456_),
    .B(_2457_),
    .CIN(_2458_),
    .COUT(_2459_),
    .SUM(_2460_));
 sky130_fd_sc_hs__fa_1 _7375_ (.A(_2461_),
    .B(_2462_),
    .CIN(_2463_),
    .COUT(_2464_),
    .SUM(_2465_));
 sky130_fd_sc_hs__fa_1 _7376_ (.A(_2466_),
    .B(_2467_),
    .CIN(_2468_),
    .COUT(_2469_),
    .SUM(_2470_));
 sky130_fd_sc_hs__fa_1 _7377_ (.A(_2470_),
    .B(_2421_),
    .CIN(_2460_),
    .COUT(_2471_),
    .SUM(_2472_));
 sky130_fd_sc_hs__fa_1 _7378_ (.A(_2473_),
    .B(_2474_),
    .CIN(_2475_),
    .COUT(_2476_),
    .SUM(_2477_));
 sky130_fd_sc_hs__fa_2 _7379_ (.A(_2478_),
    .B(_2438_),
    .CIN(_2477_),
    .COUT(_2479_),
    .SUM(_2480_));
 sky130_fd_sc_hs__fa_1 _7380_ (.A(_2481_),
    .B(_2480_),
    .CIN(_2482_),
    .COUT(_2483_),
    .SUM(_2484_));
 sky130_fd_sc_hs__fa_1 _7381_ (.A(_2485_),
    .B(_2433_),
    .CIN(_2472_),
    .COUT(_2486_),
    .SUM(_2487_));
 sky130_fd_sc_hs__fa_1 _7382_ (.A(_2488_),
    .B(_2441_),
    .CIN(_2487_),
    .COUT(_2489_),
    .SUM(_2490_));
 sky130_fd_sc_hs__fa_1 _7383_ (.A(_2491_),
    .B(_2492_),
    .CIN(_2493_),
    .COUT(_2494_),
    .SUM(_2495_));
 sky130_fd_sc_hs__fa_1 _7384_ (.A(_2496_),
    .B(_2497_),
    .CIN(_2498_),
    .COUT(_2499_),
    .SUM(_2500_));
 sky130_fd_sc_hs__fa_1 _7385_ (.A(_2501_),
    .B(_2502_),
    .CIN(_2503_),
    .COUT(_2504_),
    .SUM(_2505_));
 sky130_fd_sc_hs__fa_1 _7386_ (.A(_2506_),
    .B(_2507_),
    .CIN(_2508_),
    .COUT(_2509_),
    .SUM(_2510_));
 sky130_fd_sc_hs__fa_1 _7387_ (.A(_2511_),
    .B(_2512_),
    .CIN(_2513_),
    .COUT(_2514_),
    .SUM(_2515_));
 sky130_fd_sc_hs__fa_1 _7388_ (.A(_2515_),
    .B(_2459_),
    .CIN(_2505_),
    .COUT(_2516_),
    .SUM(_2517_));
 sky130_fd_sc_hs__fa_1 _7389_ (.A(_2518_),
    .B(_2519_),
    .CIN(_2520_),
    .COUT(_2521_),
    .SUM(_2522_));
 sky130_fd_sc_hs__fa_2 _7390_ (.A(_2523_),
    .B(_2524_),
    .CIN(_2525_),
    .COUT(_2526_),
    .SUM(_2527_));
 sky130_fd_sc_hs__fa_1 _7391_ (.A(_2528_),
    .B(_2527_),
    .CIN(_2469_),
    .COUT(_2529_),
    .SUM(_2530_));
 sky130_fd_sc_hs__fa_1 _7392_ (.A(_2530_),
    .B(_2471_),
    .CIN(_2517_),
    .COUT(_2531_),
    .SUM(_2532_));
 sky130_fd_sc_hs__fa_1 _7393_ (.A(_2483_),
    .B(_2533_),
    .CIN(_2534_),
    .COUT(_2535_),
    .SUM(_2536_));
 sky130_fd_sc_hs__fa_1 _7394_ (.A(_2537_),
    .B(_2538_),
    .CIN(_2539_),
    .COUT(_2540_),
    .SUM(_2541_));
 sky130_fd_sc_hs__fa_1 _7395_ (.A(_2542_),
    .B(_2543_),
    .CIN(_2544_),
    .COUT(_2545_),
    .SUM(_2546_));
 sky130_fd_sc_hs__fa_1 _7396_ (.A(_2547_),
    .B(_2548_),
    .CIN(_2549_),
    .COUT(_2550_),
    .SUM(_2551_));
 sky130_fd_sc_hs__fa_1 _7397_ (.A(_2552_),
    .B(_2553_),
    .CIN(_2554_),
    .COUT(_2555_),
    .SUM(_2556_));
 sky130_fd_sc_hs__fa_2 _7398_ (.A(_2557_),
    .B(_2558_),
    .CIN(_2559_),
    .COUT(_2560_),
    .SUM(_2561_));
 sky130_fd_sc_hs__fa_1 _7399_ (.A(_2561_),
    .B(_2504_),
    .CIN(_2551_),
    .COUT(_2562_),
    .SUM(_2563_));
 sky130_fd_sc_hs__fa_1 _7400_ (.A(_2564_),
    .B(_2565_),
    .CIN(_2566_),
    .COUT(_2567_),
    .SUM(_2568_));
 sky130_fd_sc_hs__fa_1 _7401_ (.A(_2569_),
    .B(_2570_),
    .CIN(_2571_),
    .COUT(_2572_),
    .SUM(_2573_));
 sky130_fd_sc_hs__fa_1 _7402_ (.A(_2574_),
    .B(_2575_),
    .CIN(_2576_),
    .COUT(_2577_),
    .SUM(_2578_));
 sky130_fd_sc_hs__fa_1 _7403_ (.A(_2579_),
    .B(_2580_),
    .CIN(_2581_),
    .COUT(_2582_),
    .SUM(_2583_));
 sky130_fd_sc_hs__fa_1 _7404_ (.A(_2584_),
    .B(_2516_),
    .CIN(_2563_),
    .COUT(_2585_),
    .SUM(_2586_));
 sky130_fd_sc_hs__fa_1 _7405_ (.A(_2587_),
    .B(_2588_),
    .CIN(_2589_),
    .COUT(_2590_),
    .SUM(_2591_));
 sky130_fd_sc_hs__fa_1 _7406_ (.A(_2592_),
    .B(_2593_),
    .CIN(_2594_),
    .COUT(_2595_),
    .SUM(_2596_));
 sky130_fd_sc_hs__fa_1 _7407_ (.A(_2597_),
    .B(_2598_),
    .CIN(_2599_),
    .COUT(_2600_),
    .SUM(_2601_));
 sky130_fd_sc_hs__fa_1 _7408_ (.A(_2602_),
    .B(_2603_),
    .CIN(_2604_),
    .COUT(_2605_),
    .SUM(_2606_));
 sky130_fd_sc_hs__fa_1 _7409_ (.A(_2607_),
    .B(_2608_),
    .CIN(_2609_),
    .COUT(_2610_),
    .SUM(_2611_));
 sky130_fd_sc_hs__fa_2 _7410_ (.A(_2612_),
    .B(_2613_),
    .CIN(_2614_),
    .COUT(_2615_),
    .SUM(_2616_));
 sky130_fd_sc_hs__fa_1 _7411_ (.A(_2616_),
    .B(_2550_),
    .CIN(_2606_),
    .COUT(_2617_),
    .SUM(_2618_));
 sky130_fd_sc_hs__fa_1 _7412_ (.A(_2619_),
    .B(_2620_),
    .CIN(_2621_),
    .COUT(_2622_),
    .SUM(_2623_));
 sky130_fd_sc_hs__fa_1 _7413_ (.A(_2624_),
    .B(_2625_),
    .CIN(_2626_),
    .COUT(_2627_),
    .SUM(_2628_));
 sky130_fd_sc_hs__fa_1 _7414_ (.A(_2629_),
    .B(_2630_),
    .CIN(_2631_),
    .COUT(_2632_),
    .SUM(_2633_));
 sky130_fd_sc_hs__fa_1 _7415_ (.A(_2634_),
    .B(_2635_),
    .CIN(_2636_),
    .COUT(_2637_),
    .SUM(_2638_));
 sky130_fd_sc_hs__fa_1 _7416_ (.A(_2639_),
    .B(_2562_),
    .CIN(_2618_),
    .COUT(_2640_),
    .SUM(_2641_));
 sky130_fd_sc_hs__fa_1 _7417_ (.A(_2642_),
    .B(_2585_),
    .CIN(_2641_),
    .COUT(_2643_),
    .SUM(_2644_));
 sky130_fd_sc_hs__fa_1 _7418_ (.A(_2645_),
    .B(_2646_),
    .CIN(_2644_),
    .COUT(_2647_),
    .SUM(_2648_));
 sky130_fd_sc_hs__fa_1 _7419_ (.A(_2650_),
    .B(_2651_),
    .CIN(_2652_),
    .COUT(_2653_),
    .SUM(_2654_));
 sky130_fd_sc_hs__fa_1 _7420_ (.A(_2655_),
    .B(_2656_),
    .CIN(_2657_),
    .COUT(_2658_),
    .SUM(_2659_));
 sky130_fd_sc_hs__fa_1 _7421_ (.A(_2660_),
    .B(_2661_),
    .CIN(_2662_),
    .COUT(_2663_),
    .SUM(_2664_));
 sky130_fd_sc_hs__fa_1 _7422_ (.A(_2665_),
    .B(_2666_),
    .CIN(_2667_),
    .COUT(_2668_),
    .SUM(_2669_));
 sky130_fd_sc_hs__fa_1 _7423_ (.A(_2670_),
    .B(_2671_),
    .CIN(_2672_),
    .COUT(_2673_),
    .SUM(_2674_));
 sky130_fd_sc_hs__fa_1 _7424_ (.A(_2674_),
    .B(_2605_),
    .CIN(_2664_),
    .COUT(_2675_),
    .SUM(_2676_));
 sky130_fd_sc_hs__fa_1 _7425_ (.A(_2677_),
    .B(_2678_),
    .CIN(_2679_),
    .COUT(_2680_),
    .SUM(_2681_));
 sky130_fd_sc_hs__fa_1 _7426_ (.A(_2682_),
    .B(_2683_),
    .CIN(_2684_),
    .COUT(_2685_),
    .SUM(_2686_));
 sky130_fd_sc_hs__fa_1 _7427_ (.A(_2687_),
    .B(_2688_),
    .CIN(_2689_),
    .COUT(_2690_),
    .SUM(_2691_));
 sky130_fd_sc_hs__fa_2 _7428_ (.A(_2632_),
    .B(_2691_),
    .CIN(_2615_),
    .COUT(_2692_),
    .SUM(_2693_));
 sky130_fd_sc_hs__fa_1 _7429_ (.A(_2693_),
    .B(_2617_),
    .CIN(_2676_),
    .COUT(_2694_),
    .SUM(_2695_));
 sky130_fd_sc_hs__fa_1 _7430_ (.A(_2696_),
    .B(_2640_),
    .CIN(_2695_),
    .COUT(_2697_),
    .SUM(_2698_));
 sky130_fd_sc_hs__fa_1 _7431_ (.A(_2699_),
    .B(_2643_),
    .CIN(_2698_),
    .COUT(_2700_),
    .SUM(_2701_));
 sky130_fd_sc_hs__fa_1 _7432_ (.A(_2703_),
    .B(_2704_),
    .CIN(_2705_),
    .COUT(_2706_),
    .SUM(_2707_));
 sky130_fd_sc_hs__fa_1 _7433_ (.A(_2708_),
    .B(_2709_),
    .CIN(_2710_),
    .COUT(_2711_),
    .SUM(_2712_));
 sky130_fd_sc_hs__fa_1 _7434_ (.A(_2713_),
    .B(_2714_),
    .CIN(_2715_),
    .COUT(_2716_),
    .SUM(_2717_));
 sky130_fd_sc_hs__fa_1 _7435_ (.A(_2718_),
    .B(_2719_),
    .CIN(_2720_),
    .COUT(_2721_),
    .SUM(_2722_));
 sky130_fd_sc_hs__fa_2 _7436_ (.A(_2723_),
    .B(_2724_),
    .CIN(_2725_),
    .COUT(_2726_),
    .SUM(_2727_));
 sky130_fd_sc_hs__fa_1 _7437_ (.A(_2727_),
    .B(_2663_),
    .CIN(_2717_),
    .COUT(_2728_),
    .SUM(_2729_));
 sky130_fd_sc_hs__fa_1 _7438_ (.A(_2730_),
    .B(_2731_),
    .CIN(_2732_),
    .COUT(_2733_),
    .SUM(_2734_));
 sky130_fd_sc_hs__fa_1 _7439_ (.A(_2735_),
    .B(_2736_),
    .CIN(_2737_),
    .COUT(_2738_),
    .SUM(_2739_));
 sky130_fd_sc_hs__fa_1 _7440_ (.A(_2740_),
    .B(_2741_),
    .CIN(_2742_),
    .COUT(_2743_),
    .SUM(_2744_));
 sky130_fd_sc_hs__fa_1 _7441_ (.A(_2690_),
    .B(_2744_),
    .CIN(_2673_),
    .COUT(_2745_),
    .SUM(_2746_));
 sky130_fd_sc_hs__fa_1 _7442_ (.A(_2746_),
    .B(_2675_),
    .CIN(_2729_),
    .COUT(_2747_),
    .SUM(_2748_));
 sky130_fd_sc_hs__fa_1 _7443_ (.A(_2749_),
    .B(_2750_),
    .CIN(_2751_),
    .COUT(_2752_),
    .SUM(_2753_));
 sky130_fd_sc_hs__fa_1 _7444_ (.A(_2754_),
    .B(_2753_),
    .CIN(_2685_),
    .COUT(_2755_),
    .SUM(_2756_));
 sky130_fd_sc_hs__fa_1 _7445_ (.A(_2757_),
    .B(_2758_),
    .CIN(_2759_),
    .COUT(_2760_),
    .SUM(_2761_));
 sky130_fd_sc_hs__fa_1 _7446_ (.A(_2762_),
    .B(_2763_),
    .CIN(_2764_),
    .COUT(_2765_),
    .SUM(_2766_));
 sky130_fd_sc_hs__fa_1 _7447_ (.A(_2767_),
    .B(_2694_),
    .CIN(_2748_),
    .COUT(_2768_),
    .SUM(_2769_));
 sky130_fd_sc_hs__fa_2 _7448_ (.A(_2770_),
    .B(_2697_),
    .CIN(_2769_),
    .COUT(_2771_),
    .SUM(_2772_));
 sky130_fd_sc_hs__fa_1 _7449_ (.A(_2774_),
    .B(_2775_),
    .CIN(_2703_),
    .COUT(_2776_),
    .SUM(_2777_));
 sky130_fd_sc_hs__fa_1 _7450_ (.A(_2780_),
    .B(_2781_),
    .CIN(_2782_),
    .COUT(_2783_),
    .SUM(_2784_));
 sky130_fd_sc_hs__fa_1 _7451_ (.A(_2785_),
    .B(_2786_),
    .CIN(_2787_),
    .COUT(_2788_),
    .SUM(_2789_));
 sky130_fd_sc_hs__fa_1 _7452_ (.A(_2790_),
    .B(_2791_),
    .CIN(_2792_),
    .COUT(_2793_),
    .SUM(_2794_));
 sky130_fd_sc_hs__fa_2 _7453_ (.A(_2795_),
    .B(_2796_),
    .CIN(_2797_),
    .COUT(_2798_),
    .SUM(_2799_));
 sky130_fd_sc_hs__fa_1 _7454_ (.A(_2799_),
    .B(_2716_),
    .CIN(_2789_),
    .COUT(_2800_),
    .SUM(_2801_));
 sky130_fd_sc_hs__fa_1 _7455_ (.A(_2802_),
    .B(_2803_),
    .CIN(_2804_),
    .COUT(_2805_),
    .SUM(_2806_));
 sky130_fd_sc_hs__fa_1 _7456_ (.A(_2807_),
    .B(_2808_),
    .CIN(_2809_),
    .COUT(_2810_),
    .SUM(_2811_));
 sky130_fd_sc_hs__fa_1 _7457_ (.A(_2812_),
    .B(_2813_),
    .CIN(_2814_),
    .COUT(_2815_),
    .SUM(_2816_));
 sky130_fd_sc_hs__fa_2 _7458_ (.A(_2743_),
    .B(_2816_),
    .CIN(_2726_),
    .COUT(_2817_),
    .SUM(_2818_));
 sky130_fd_sc_hs__fa_1 _7459_ (.A(_2818_),
    .B(_2728_),
    .CIN(_2801_),
    .COUT(_2819_),
    .SUM(_2820_));
 sky130_fd_sc_hs__fa_1 _7460_ (.A(_2821_),
    .B(_2822_),
    .CIN(_2823_),
    .COUT(_2824_),
    .SUM(_2825_));
 sky130_fd_sc_hs__fa_1 _7461_ (.A(_2826_),
    .B(_2827_),
    .CIN(_2828_),
    .COUT(_2829_),
    .SUM(_2830_));
 sky130_fd_sc_hs__fa_1 _7462_ (.A(_2760_),
    .B(_2831_),
    .CIN(_2745_),
    .COUT(_2832_),
    .SUM(_2833_));
 sky130_fd_sc_hs__fa_1 _7463_ (.A(_2833_),
    .B(_2747_),
    .CIN(_2820_),
    .COUT(_2834_),
    .SUM(_2835_));
 sky130_fd_sc_hs__fa_2 _7464_ (.A(_2836_),
    .B(_2768_),
    .CIN(_2835_),
    .COUT(_2837_),
    .SUM(_2838_));
 sky130_fd_sc_hs__fa_1 _7465_ (.A(_2839_),
    .B(_2774_),
    .CIN(_2703_),
    .COUT(_2840_),
    .SUM(_2841_));
 sky130_fd_sc_hs__fa_1 _7466_ (.A(_2842_),
    .B(_2843_),
    .CIN(_2844_),
    .COUT(_2845_),
    .SUM(_2846_));
 sky130_fd_sc_hs__fa_1 _7467_ (.A(_2847_),
    .B(_2848_),
    .CIN(_2849_),
    .COUT(_2850_),
    .SUM(_2851_));
 sky130_fd_sc_hs__fa_1 _7468_ (.A(_2852_),
    .B(_2853_),
    .CIN(_2854_),
    .COUT(_2855_),
    .SUM(_2856_));
 sky130_fd_sc_hs__fa_1 _7469_ (.A(_2857_),
    .B(_2858_),
    .CIN(_2859_),
    .COUT(_2860_),
    .SUM(_2861_));
 sky130_fd_sc_hs__fa_1 _7470_ (.A(_2861_),
    .B(_2788_),
    .CIN(_2851_),
    .COUT(_2862_),
    .SUM(_2863_));
 sky130_fd_sc_hs__fa_1 _7471_ (.A(_2864_),
    .B(_2865_),
    .CIN(_2866_),
    .COUT(_2867_),
    .SUM(_2868_));
 sky130_fd_sc_hs__fa_1 _7472_ (.A(_2869_),
    .B(_2870_),
    .CIN(_2871_),
    .COUT(_2872_),
    .SUM(_2873_));
 sky130_fd_sc_hs__fa_1 _7473_ (.A(_2874_),
    .B(_2875_),
    .CIN(_2876_),
    .COUT(_2877_),
    .SUM(_2878_));
 sky130_fd_sc_hs__fa_1 _7474_ (.A(_2815_),
    .B(_2878_),
    .CIN(_2798_),
    .COUT(_2879_),
    .SUM(_2880_));
 sky130_fd_sc_hs__fa_1 _7475_ (.A(_2880_),
    .B(_2800_),
    .CIN(_2863_),
    .COUT(_2881_),
    .SUM(_2882_));
 sky130_fd_sc_hs__fa_1 _7476_ (.A(_2883_),
    .B(_2884_),
    .CIN(_2885_),
    .COUT(_2886_),
    .SUM(_2887_));
 sky130_fd_sc_hs__fa_1 _7477_ (.A(_2888_),
    .B(_2889_),
    .CIN(_2890_),
    .COUT(_2891_),
    .SUM(_2892_));
 sky130_fd_sc_hs__fa_1 _7478_ (.A(_2893_),
    .B(_2894_),
    .CIN(_2895_),
    .COUT(_2896_),
    .SUM(_2897_));
 sky130_fd_sc_hs__fa_1 _7479_ (.A(_2898_),
    .B(_2819_),
    .CIN(_2882_),
    .COUT(_2899_),
    .SUM(_2900_));
 sky130_fd_sc_hs__fa_1 _7480_ (.A(_2832_),
    .B(_2834_),
    .CIN(_2900_),
    .COUT(_2901_),
    .SUM(_2902_));
 sky130_fd_sc_hs__fa_1 _7481_ (.A(_2903_),
    .B(_2774_),
    .CIN(_2703_),
    .COUT(_2904_),
    .SUM(_2905_));
 sky130_fd_sc_hs__fa_1 _7482_ (.A(_2906_),
    .B(_2907_),
    .CIN(_2844_),
    .COUT(_2908_),
    .SUM(_2909_));
 sky130_fd_sc_hs__fa_1 _7483_ (.A(_2910_),
    .B(_2911_),
    .CIN(_2912_),
    .COUT(_2913_),
    .SUM(_2914_));
 sky130_fd_sc_hs__fa_1 _7484_ (.A(_2915_),
    .B(_2916_),
    .CIN(_2917_),
    .COUT(_2918_),
    .SUM(_2919_));
 sky130_fd_sc_hs__fa_1 _7485_ (.A(_2920_),
    .B(_2921_),
    .CIN(_2922_),
    .COUT(_2923_),
    .SUM(_2924_));
 sky130_fd_sc_hs__fa_1 _7486_ (.A(_2924_),
    .B(_2850_),
    .CIN(_2914_),
    .COUT(_2925_),
    .SUM(_2926_));
 sky130_fd_sc_hs__fa_1 _7487_ (.A(_2927_),
    .B(_2928_),
    .CIN(_2929_),
    .COUT(_2930_),
    .SUM(_2931_));
 sky130_fd_sc_hs__fa_1 _7488_ (.A(_2932_),
    .B(_2933_),
    .CIN(_2934_),
    .COUT(_2935_),
    .SUM(_2936_));
 sky130_fd_sc_hs__fa_1 _7489_ (.A(_2937_),
    .B(_2938_),
    .CIN(_2939_),
    .COUT(_2940_),
    .SUM(_2941_));
 sky130_fd_sc_hs__fa_2 _7490_ (.A(_2877_),
    .B(_2941_),
    .CIN(_2860_),
    .COUT(_2942_),
    .SUM(_2943_));
 sky130_fd_sc_hs__fa_2 _7491_ (.A(_2943_),
    .B(_2862_),
    .CIN(_2926_),
    .COUT(_2944_),
    .SUM(_2945_));
 sky130_fd_sc_hs__fa_1 _7492_ (.A(_2946_),
    .B(_2947_),
    .CIN(_2948_),
    .COUT(_2949_),
    .SUM(_2950_));
 sky130_fd_sc_hs__fa_1 _7493_ (.A(_2951_),
    .B(_2952_),
    .CIN(_2953_),
    .COUT(_2954_),
    .SUM(_2955_));
 sky130_fd_sc_hs__fa_1 _7494_ (.A(_2956_),
    .B(_2957_),
    .CIN(_2958_),
    .COUT(_2959_),
    .SUM(_2960_));
 sky130_fd_sc_hs__fa_2 _7495_ (.A(_2961_),
    .B(_2881_),
    .CIN(_2945_),
    .COUT(_2962_),
    .SUM(_2963_));
 sky130_fd_sc_hs__fa_2 _7496_ (.A(_2964_),
    .B(_2899_),
    .CIN(_2963_),
    .COUT(_2965_),
    .SUM(_2966_));
 sky130_fd_sc_hs__fa_1 _7497_ (.A(_2967_),
    .B(_2774_),
    .CIN(_2703_),
    .COUT(_2968_),
    .SUM(_2969_));
 sky130_fd_sc_hs__fa_4 _7498_ (.A(_2970_),
    .B(_2907_),
    .CIN(_2844_),
    .COUT(_2971_),
    .SUM(_2972_));
 sky130_fd_sc_hs__fa_1 _7499_ (.A(_2973_),
    .B(_2974_),
    .CIN(_2975_),
    .COUT(_2976_),
    .SUM(_2977_));
 sky130_fd_sc_hs__fa_1 _7500_ (.A(_2978_),
    .B(_2979_),
    .CIN(_2980_),
    .COUT(_2981_),
    .SUM(_2982_));
 sky130_fd_sc_hs__fa_2 _7501_ (.A(_2983_),
    .B(_2984_),
    .CIN(_2985_),
    .COUT(_2986_),
    .SUM(_2987_));
 sky130_fd_sc_hs__fa_1 _7502_ (.A(_2987_),
    .B(_2913_),
    .CIN(_2977_),
    .COUT(_2988_),
    .SUM(_2989_));
 sky130_fd_sc_hs__fa_1 _7503_ (.A(_2990_),
    .B(_2991_),
    .CIN(_2992_),
    .COUT(_2993_),
    .SUM(_2994_));
 sky130_fd_sc_hs__fa_1 _7504_ (.A(_2995_),
    .B(_2996_),
    .CIN(_2997_),
    .COUT(_2998_),
    .SUM(_2999_));
 sky130_fd_sc_hs__fa_1 _7505_ (.A(_3000_),
    .B(_3001_),
    .CIN(_3002_),
    .COUT(_3003_),
    .SUM(_3004_));
 sky130_fd_sc_hs__fa_2 _7506_ (.A(_2940_),
    .B(_3004_),
    .CIN(_2923_),
    .COUT(_3005_),
    .SUM(_3006_));
 sky130_fd_sc_hs__fa_1 _7507_ (.A(_3006_),
    .B(_2925_),
    .CIN(_2989_),
    .COUT(_3007_),
    .SUM(_3008_));
 sky130_fd_sc_hs__fa_1 _7508_ (.A(_3009_),
    .B(_3010_),
    .CIN(_3011_),
    .COUT(_3012_),
    .SUM(_3013_));
 sky130_fd_sc_hs__fa_1 _7509_ (.A(_3014_),
    .B(_3015_),
    .CIN(_3016_),
    .COUT(_3017_),
    .SUM(_3018_));
 sky130_fd_sc_hs__fa_1 _7510_ (.A(_3019_),
    .B(_3020_),
    .CIN(_3021_),
    .COUT(_3022_),
    .SUM(_3023_));
 sky130_fd_sc_hs__fa_1 _7511_ (.A(_3024_),
    .B(_2944_),
    .CIN(_3008_),
    .COUT(_3025_),
    .SUM(_3026_));
 sky130_fd_sc_hs__fa_1 _7512_ (.A(_3027_),
    .B(_2962_),
    .CIN(_3026_),
    .COUT(_3028_),
    .SUM(_3029_));
 sky130_fd_sc_hs__fa_1 _7513_ (.A(_3030_),
    .B(_2774_),
    .CIN(_2703_),
    .COUT(_3031_),
    .SUM(_3032_));
 sky130_fd_sc_hs__fa_1 _7514_ (.A(_3033_),
    .B(_3034_),
    .CIN(_2973_),
    .COUT(_3035_),
    .SUM(_3036_));
 sky130_fd_sc_hs__fa_1 _7515_ (.A(_3037_),
    .B(_3038_),
    .CIN(_3039_),
    .COUT(_3040_),
    .SUM(_3041_));
 sky130_fd_sc_hs__fa_2 _7516_ (.A(_3042_),
    .B(_3043_),
    .CIN(_3044_),
    .COUT(_3045_),
    .SUM(_3046_));
 sky130_fd_sc_hs__fa_1 _7517_ (.A(_3046_),
    .B(_2976_),
    .CIN(_3036_),
    .COUT(_3047_),
    .SUM(_3048_));
 sky130_fd_sc_hs__fa_1 _7518_ (.A(_3049_),
    .B(_3050_),
    .CIN(_3051_),
    .COUT(_3052_),
    .SUM(_3053_));
 sky130_fd_sc_hs__fa_1 _7519_ (.A(_3054_),
    .B(_3055_),
    .CIN(_3056_),
    .COUT(_3057_),
    .SUM(_3058_));
 sky130_fd_sc_hs__fa_1 _7520_ (.A(_3059_),
    .B(_3060_),
    .CIN(_3061_),
    .COUT(_3062_),
    .SUM(_3063_));
 sky130_fd_sc_hs__fa_2 _7521_ (.A(_3003_),
    .B(_3063_),
    .CIN(_2986_),
    .COUT(_3064_),
    .SUM(_3065_));
 sky130_fd_sc_hs__fa_1 _7522_ (.A(_3065_),
    .B(_2988_),
    .CIN(_3048_),
    .COUT(_3066_),
    .SUM(_3067_));
 sky130_fd_sc_hs__fa_1 _7523_ (.A(_3068_),
    .B(_3069_),
    .CIN(_3070_),
    .COUT(_3071_),
    .SUM(_3072_));
 sky130_fd_sc_hs__fa_1 _7524_ (.A(_3073_),
    .B(_3074_),
    .CIN(_3075_),
    .COUT(_3076_),
    .SUM(_3077_));
 sky130_fd_sc_hs__fa_1 _7525_ (.A(_3078_),
    .B(_3079_),
    .CIN(_3080_),
    .COUT(_3081_),
    .SUM(_3082_));
 sky130_fd_sc_hs__fa_1 _7526_ (.A(_3083_),
    .B(_3007_),
    .CIN(_3067_),
    .COUT(_3084_),
    .SUM(_3085_));
 sky130_fd_sc_hs__fa_1 _7527_ (.A(_3086_),
    .B(_3025_),
    .CIN(_3085_),
    .COUT(_3087_),
    .SUM(_3088_));
 sky130_fd_sc_hs__fa_1 _7528_ (.A(_3089_),
    .B(_2778_),
    .CIN(_2779_),
    .COUT(_3090_),
    .SUM(_3091_));
 sky130_fd_sc_hs__fa_1 _7529_ (.A(_3031_),
    .B(_3092_),
    .CIN(_2972_),
    .COUT(_3093_),
    .SUM(_3094_));
 sky130_fd_sc_hs__fa_1 _7530_ (.A(_3095_),
    .B(_3096_),
    .CIN(_3039_),
    .COUT(_3097_),
    .SUM(_3098_));
 sky130_fd_sc_hs__fa_2 _7531_ (.A(_3099_),
    .B(_3100_),
    .CIN(_3044_),
    .COUT(_3101_),
    .SUM(_3102_));
 sky130_fd_sc_hs__fa_1 _7532_ (.A(_3102_),
    .B(_3035_),
    .CIN(_3103_),
    .COUT(_3104_),
    .SUM(_3105_));
 sky130_fd_sc_hs__fa_1 _7533_ (.A(_3106_),
    .B(_3107_),
    .CIN(_3108_),
    .COUT(_3109_),
    .SUM(_3110_));
 sky130_fd_sc_hs__fa_1 _7534_ (.A(_3111_),
    .B(_3112_),
    .CIN(_3113_),
    .COUT(_3114_),
    .SUM(_3115_));
 sky130_fd_sc_hs__fa_1 _7535_ (.A(_3116_),
    .B(_3117_),
    .CIN(_3118_),
    .COUT(_3119_),
    .SUM(_3120_));
 sky130_fd_sc_hs__fa_2 _7536_ (.A(_3062_),
    .B(_3120_),
    .CIN(_3045_),
    .COUT(_3121_),
    .SUM(_3122_));
 sky130_fd_sc_hs__fa_1 _7537_ (.A(_3122_),
    .B(_3047_),
    .CIN(_3105_),
    .COUT(_3123_),
    .SUM(_3124_));
 sky130_fd_sc_hs__fa_1 _7538_ (.A(_3125_),
    .B(_3126_),
    .CIN(_3127_),
    .COUT(_3128_),
    .SUM(_3129_));
 sky130_fd_sc_hs__fa_1 _7539_ (.A(_3130_),
    .B(_3131_),
    .CIN(_3132_),
    .COUT(_3133_),
    .SUM(_3134_));
 sky130_fd_sc_hs__fa_1 _7540_ (.A(_3135_),
    .B(_3136_),
    .CIN(_3137_),
    .COUT(_3138_),
    .SUM(_3139_));
 sky130_fd_sc_hs__fa_1 _7541_ (.A(_3140_),
    .B(_3066_),
    .CIN(_3124_),
    .COUT(_3141_),
    .SUM(_3142_));
 sky130_fd_sc_hs__fa_1 _7542_ (.A(_3143_),
    .B(_3084_),
    .CIN(_3142_),
    .COUT(_3144_),
    .SUM(_3145_));
 sky130_fd_sc_hs__fa_1 _7543_ (.A(_3146_),
    .B(_2778_),
    .CIN(_2779_),
    .COUT(_3147_),
    .SUM(_3148_));
 sky130_fd_sc_hs__fa_1 _7544_ (.A(_3149_),
    .B(_3150_),
    .CIN(_2972_),
    .COUT(_3151_),
    .SUM(_3152_));
 sky130_fd_sc_hs__fa_1 _7545_ (.A(_3153_),
    .B(_3096_),
    .CIN(_3039_),
    .COUT(_3154_),
    .SUM(_3155_));
 sky130_fd_sc_hs__fa_1 _7546_ (.A(_3156_),
    .B(_3157_),
    .CIN(_3044_),
    .COUT(_3158_),
    .SUM(_3159_));
 sky130_fd_sc_hs__fa_1 _7547_ (.A(_3159_),
    .B(_3160_),
    .CIN(_3161_),
    .COUT(_3162_),
    .SUM(_3163_));
 sky130_fd_sc_hs__fa_1 _7548_ (.A(_3164_),
    .B(_3165_),
    .CIN(_3166_),
    .COUT(_3167_),
    .SUM(_3168_));
 sky130_fd_sc_hs__fa_1 _7549_ (.A(_3169_),
    .B(_3170_),
    .CIN(_3171_),
    .COUT(_3172_),
    .SUM(_3173_));
 sky130_fd_sc_hs__fa_1 _7550_ (.A(_3174_),
    .B(_3175_),
    .CIN(_3176_),
    .COUT(_3177_),
    .SUM(_3178_));
 sky130_fd_sc_hs__fa_2 _7551_ (.A(_3119_),
    .B(_3178_),
    .CIN(_3101_),
    .COUT(_3179_),
    .SUM(_3180_));
 sky130_fd_sc_hs__fa_1 _7552_ (.A(_3180_),
    .B(_3104_),
    .CIN(_3163_),
    .COUT(_3181_),
    .SUM(_3182_));
 sky130_fd_sc_hs__fa_1 _7553_ (.A(_3183_),
    .B(_3184_),
    .CIN(_3185_),
    .COUT(_3186_),
    .SUM(_3187_));
 sky130_fd_sc_hs__fa_1 _7554_ (.A(_3188_),
    .B(_3189_),
    .CIN(_3190_),
    .COUT(_3191_),
    .SUM(_3192_));
 sky130_fd_sc_hs__fa_1 _7555_ (.A(_3193_),
    .B(_3194_),
    .CIN(_3195_),
    .COUT(_3196_),
    .SUM(_3197_));
 sky130_fd_sc_hs__fa_1 _7556_ (.A(_3198_),
    .B(_3123_),
    .CIN(_3182_),
    .COUT(_3199_),
    .SUM(_3200_));
 sky130_fd_sc_hs__fa_1 _7557_ (.A(_3201_),
    .B(_3141_),
    .CIN(_3200_),
    .COUT(_3202_),
    .SUM(_3203_));
 sky130_fd_sc_hs__fa_1 _7558_ (.A(_3204_),
    .B(_2778_),
    .CIN(_2779_),
    .COUT(_3205_),
    .SUM(_3206_));
 sky130_fd_sc_hs__fa_1 _7559_ (.A(_3207_),
    .B(_3208_),
    .CIN(_2972_),
    .COUT(_3209_),
    .SUM(_3210_));
 sky130_fd_sc_hs__fa_4 _7560_ (.A(_3211_),
    .B(_3157_),
    .CIN(_3044_),
    .COUT(_3212_),
    .SUM(_3213_));
 sky130_fd_sc_hs__fa_1 _7561_ (.A(_3213_),
    .B(_3214_),
    .CIN(_3215_),
    .COUT(_3216_),
    .SUM(_3217_));
 sky130_fd_sc_hs__fa_1 _7562_ (.A(_3218_),
    .B(_3219_),
    .CIN(_3220_),
    .COUT(_3221_),
    .SUM(_3222_));
 sky130_fd_sc_hs__fa_1 _7563_ (.A(_3223_),
    .B(_3224_),
    .CIN(_3225_),
    .COUT(_3226_),
    .SUM(_3227_));
 sky130_fd_sc_hs__fa_1 _7564_ (.A(_3228_),
    .B(_3229_),
    .CIN(_3230_),
    .COUT(_3231_),
    .SUM(_3232_));
 sky130_fd_sc_hs__fa_2 _7565_ (.A(_3177_),
    .B(_3232_),
    .CIN(_3158_),
    .COUT(_3233_),
    .SUM(_3234_));
 sky130_fd_sc_hs__fa_1 _7566_ (.A(_3234_),
    .B(_3162_),
    .CIN(_3217_),
    .COUT(_3235_),
    .SUM(_3236_));
 sky130_fd_sc_hs__fa_1 _7567_ (.A(_3237_),
    .B(_3238_),
    .CIN(_3239_),
    .COUT(_3240_),
    .SUM(_3241_));
 sky130_fd_sc_hs__fa_1 _7568_ (.A(_3242_),
    .B(_3243_),
    .CIN(_3244_),
    .COUT(_3245_),
    .SUM(_3246_));
 sky130_fd_sc_hs__fa_1 _7569_ (.A(_3247_),
    .B(_3248_),
    .CIN(_3249_),
    .COUT(_3250_),
    .SUM(_3251_));
 sky130_fd_sc_hs__fa_1 _7570_ (.A(_3252_),
    .B(_3181_),
    .CIN(_3236_),
    .COUT(_3253_),
    .SUM(_3254_));
 sky130_fd_sc_hs__fa_1 _7571_ (.A(_3255_),
    .B(_3199_),
    .CIN(_3254_),
    .COUT(_3256_),
    .SUM(_3257_));
 sky130_fd_sc_hs__fa_1 _7572_ (.A(_3258_),
    .B(_2774_),
    .CIN(_2703_),
    .COUT(_3259_),
    .SUM(_3260_));
 sky130_fd_sc_hs__fa_1 _7573_ (.A(_3205_),
    .B(_3261_),
    .CIN(_2973_),
    .COUT(_3262_),
    .SUM(_3263_));
 sky130_fd_sc_hs__fa_1 _7574_ (.A(_3209_),
    .B(_3264_),
    .CIN(_3265_),
    .COUT(_3266_),
    .SUM(_3267_));
 sky130_fd_sc_hs__fa_1 _7575_ (.A(_3268_),
    .B(_3269_),
    .CIN(_3220_),
    .COUT(_3270_),
    .SUM(_3271_));
 sky130_fd_sc_hs__fa_1 _7576_ (.A(_3272_),
    .B(_3273_),
    .CIN(_3274_),
    .COUT(_3275_),
    .SUM(_3276_));
 sky130_fd_sc_hs__fa_1 _7577_ (.A(_3277_),
    .B(_3278_),
    .CIN(_3279_),
    .COUT(_3280_),
    .SUM(_3281_));
 sky130_fd_sc_hs__fa_2 _7578_ (.A(_3231_),
    .B(_3281_),
    .CIN(_3212_),
    .COUT(_3282_),
    .SUM(_3283_));
 sky130_fd_sc_hs__fa_1 _7579_ (.A(_3283_),
    .B(_3216_),
    .CIN(_3284_),
    .COUT(_3285_),
    .SUM(_3286_));
 sky130_fd_sc_hs__fa_1 _7580_ (.A(_3287_),
    .B(_3288_),
    .CIN(_3289_),
    .COUT(_3290_),
    .SUM(_3291_));
 sky130_fd_sc_hs__fa_1 _7581_ (.A(_3292_),
    .B(_3293_),
    .CIN(_3294_),
    .COUT(_3295_),
    .SUM(_3296_));
 sky130_fd_sc_hs__fa_1 _7582_ (.A(_3297_),
    .B(_3298_),
    .CIN(_3299_),
    .COUT(_3300_),
    .SUM(_3301_));
 sky130_fd_sc_hs__fa_1 _7583_ (.A(_3302_),
    .B(_3235_),
    .CIN(_3286_),
    .COUT(_3303_),
    .SUM(_3304_));
 sky130_fd_sc_hs__fa_1 _7584_ (.A(_3305_),
    .B(_3253_),
    .CIN(_3304_),
    .COUT(_3306_),
    .SUM(_3307_));
 sky130_fd_sc_hs__fa_1 _7585_ (.A(_3308_),
    .B(_2778_),
    .CIN(_2779_),
    .COUT(_3309_),
    .SUM(_3310_));
 sky130_fd_sc_hs__fa_1 _7586_ (.A(_3259_),
    .B(_3311_),
    .CIN(_2972_),
    .COUT(_3312_),
    .SUM(_3313_));
 sky130_fd_sc_hs__fa_1 _7587_ (.A(_3314_),
    .B(_3313_),
    .CIN(_3265_),
    .COUT(_3315_),
    .SUM(_3316_));
 sky130_fd_sc_hs__fa_1 _7588_ (.A(_3317_),
    .B(_3269_),
    .CIN(_3220_),
    .COUT(_3318_),
    .SUM(_3319_));
 sky130_fd_sc_hs__fa_1 _7589_ (.A(_3320_),
    .B(_3321_),
    .CIN(_3322_),
    .COUT(_3323_),
    .SUM(_3324_));
 sky130_fd_sc_hs__fa_1 _7590_ (.A(_3325_),
    .B(_3326_),
    .CIN(_3327_),
    .COUT(_3328_),
    .SUM(_3329_));
 sky130_fd_sc_hs__fa_2 _7591_ (.A(_3280_),
    .B(_3329_),
    .CIN(_3212_),
    .COUT(_3330_),
    .SUM(_3331_));
 sky130_fd_sc_hs__fa_1 _7592_ (.A(_3331_),
    .B(_3332_),
    .CIN(_3333_),
    .COUT(_3334_),
    .SUM(_3335_));
 sky130_fd_sc_hs__fa_1 _7593_ (.A(_3336_),
    .B(_3337_),
    .CIN(_3338_),
    .COUT(_3339_),
    .SUM(_3340_));
 sky130_fd_sc_hs__fa_1 _7594_ (.A(_3341_),
    .B(_3342_),
    .CIN(_3343_),
    .COUT(_3344_),
    .SUM(_3345_));
 sky130_fd_sc_hs__fa_1 _7595_ (.A(_3346_),
    .B(_3347_),
    .CIN(_3348_),
    .COUT(_3349_),
    .SUM(_3350_));
 sky130_fd_sc_hs__fa_1 _7596_ (.A(_3351_),
    .B(_3285_),
    .CIN(_3335_),
    .COUT(_3352_),
    .SUM(_3353_));
 sky130_fd_sc_hs__fa_1 _7597_ (.A(_3354_),
    .B(_3303_),
    .CIN(_3353_),
    .COUT(_3355_),
    .SUM(_3356_));
 sky130_fd_sc_hs__fa_1 _7598_ (.A(_3357_),
    .B(_2778_),
    .CIN(_2779_),
    .COUT(_3358_),
    .SUM(_3359_));
 sky130_fd_sc_hs__fa_1 _7599_ (.A(_3309_),
    .B(_3359_),
    .CIN(_2973_),
    .COUT(_3360_),
    .SUM(_3361_));
 sky130_fd_sc_hs__fa_1 _7600_ (.A(_3362_),
    .B(_3361_),
    .CIN(_3213_),
    .COUT(_3363_),
    .SUM(_3364_));
 sky130_fd_sc_hs__fa_1 _7601_ (.A(_3365_),
    .B(_3366_),
    .CIN(_3367_),
    .COUT(_3368_),
    .SUM(_3369_));
 sky130_fd_sc_hs__fa_1 _7602_ (.A(_3370_),
    .B(_3371_),
    .CIN(_3327_),
    .COUT(_3372_),
    .SUM(_3373_));
 sky130_fd_sc_hs__fa_1 _7603_ (.A(_3328_),
    .B(_3373_),
    .CIN(_3212_),
    .COUT(_3374_),
    .SUM(_3375_));
 sky130_fd_sc_hs__fa_1 _7604_ (.A(_3375_),
    .B(_3376_),
    .CIN(_3364_),
    .COUT(_3377_),
    .SUM(_3378_));
 sky130_fd_sc_hs__fa_1 _7605_ (.A(_3379_),
    .B(_3380_),
    .CIN(_3381_),
    .COUT(_3382_),
    .SUM(_3383_));
 sky130_fd_sc_hs__fa_1 _7606_ (.A(_3384_),
    .B(_3385_),
    .CIN(_3386_),
    .COUT(_3387_),
    .SUM(_3388_));
 sky130_fd_sc_hs__fa_1 _7607_ (.A(_3389_),
    .B(_3390_),
    .CIN(_3391_),
    .COUT(_3392_),
    .SUM(_3393_));
 sky130_fd_sc_hs__fa_1 _7608_ (.A(_3394_),
    .B(_3334_),
    .CIN(_3378_),
    .COUT(_3395_),
    .SUM(_3396_));
 sky130_fd_sc_hs__fa_1 _7609_ (.A(_3397_),
    .B(_3352_),
    .CIN(_3396_),
    .COUT(_3398_),
    .SUM(_3399_));
 sky130_fd_sc_hs__fa_1 _7610_ (.A(_3400_),
    .B(_2778_),
    .CIN(_2779_),
    .COUT(_3401_),
    .SUM(_3402_));
 sky130_fd_sc_hs__fa_2 _7611_ (.A(_3358_),
    .B(_3402_),
    .CIN(_2973_),
    .COUT(_3403_),
    .SUM(_3404_));
 sky130_fd_sc_hs__fa_1 _7612_ (.A(_3360_),
    .B(_3404_),
    .CIN(_3213_),
    .COUT(_3405_),
    .SUM(_3406_));
 sky130_fd_sc_hs__fa_1 _7613_ (.A(_3407_),
    .B(_3408_),
    .CIN(_3367_),
    .COUT(_3409_),
    .SUM(_3410_));
 sky130_fd_sc_hs__fa_1 _7614_ (.A(_3411_),
    .B(_3371_),
    .CIN(_3327_),
    .COUT(_3412_),
    .SUM(_3413_));
 sky130_fd_sc_hs__fa_1 _7615_ (.A(_3372_),
    .B(_3413_),
    .CIN(_3212_),
    .COUT(_3414_),
    .SUM(_3415_));
 sky130_fd_sc_hs__fa_1 _7616_ (.A(_3415_),
    .B(_3363_),
    .CIN(_3406_),
    .COUT(_3416_),
    .SUM(_3417_));
 sky130_fd_sc_hs__fa_1 _7617_ (.A(_3418_),
    .B(_3419_),
    .CIN(_3420_),
    .COUT(_3421_),
    .SUM(_3422_));
 sky130_fd_sc_hs__fa_1 _7618_ (.A(_3423_),
    .B(_3424_),
    .CIN(_3425_),
    .COUT(_3426_),
    .SUM(_3427_));
 sky130_fd_sc_hs__fa_1 _7619_ (.A(_3428_),
    .B(_3429_),
    .CIN(_3430_),
    .COUT(_3431_),
    .SUM(_3432_));
 sky130_fd_sc_hs__fa_1 _7620_ (.A(_3433_),
    .B(_3377_),
    .CIN(_3417_),
    .COUT(_3434_),
    .SUM(_3435_));
 sky130_fd_sc_hs__fa_1 _7621_ (.A(_3436_),
    .B(_3395_),
    .CIN(_3435_),
    .COUT(_3437_),
    .SUM(_3438_));
 sky130_fd_sc_hs__fa_1 _7622_ (.A(_3439_),
    .B(_2778_),
    .CIN(_2779_),
    .COUT(_3440_),
    .SUM(_3441_));
 sky130_fd_sc_hs__fa_1 _7623_ (.A(_3401_),
    .B(_3441_),
    .CIN(_2973_),
    .COUT(_3442_),
    .SUM(_3443_));
 sky130_fd_sc_hs__fa_1 _7624_ (.A(_3403_),
    .B(_3443_),
    .CIN(_3213_),
    .COUT(_3444_),
    .SUM(_3445_));
 sky130_fd_sc_hs__fa_4 _7625_ (.A(_3446_),
    .B(_3408_),
    .CIN(_3367_),
    .COUT(_3447_),
    .SUM(_3448_));
 sky130_fd_sc_hs__fa_4 _7626_ (.A(_3449_),
    .B(_3371_),
    .CIN(_3327_),
    .COUT(_3450_),
    .SUM(_3451_));
 sky130_fd_sc_hs__fa_1 _7627_ (.A(_3412_),
    .B(_3451_),
    .CIN(_3212_),
    .COUT(_3452_),
    .SUM(_3453_));
 sky130_fd_sc_hs__fa_1 _7628_ (.A(_3453_),
    .B(_3405_),
    .CIN(_3445_),
    .COUT(_3454_),
    .SUM(_3455_));
 sky130_fd_sc_hs__fa_1 _7629_ (.A(_3456_),
    .B(_3457_),
    .CIN(_3458_),
    .COUT(_3459_),
    .SUM(_3460_));
 sky130_fd_sc_hs__fa_1 _7630_ (.A(_3461_),
    .B(_3462_),
    .CIN(_3463_),
    .COUT(_3464_),
    .SUM(_3465_));
 sky130_fd_sc_hs__fa_1 _7631_ (.A(_3466_),
    .B(_3467_),
    .CIN(_3468_),
    .COUT(_3469_),
    .SUM(_3470_));
 sky130_fd_sc_hs__fa_1 _7632_ (.A(_3471_),
    .B(_3416_),
    .CIN(_3455_),
    .COUT(_3472_),
    .SUM(_3473_));
 sky130_fd_sc_hs__fa_1 _7633_ (.A(_3474_),
    .B(_3434_),
    .CIN(_3473_),
    .COUT(_3475_),
    .SUM(_3476_));
 sky130_fd_sc_hs__fa_1 _7634_ (.A(_3477_),
    .B(_2778_),
    .CIN(_2779_),
    .COUT(_3478_),
    .SUM(_3479_));
 sky130_fd_sc_hs__fa_1 _7635_ (.A(_3440_),
    .B(_3479_),
    .CIN(_2973_),
    .COUT(_3480_),
    .SUM(_3481_));
 sky130_fd_sc_hs__fa_1 _7636_ (.A(_3442_),
    .B(_3481_),
    .CIN(_3213_),
    .COUT(_3482_),
    .SUM(_3483_));
 sky130_fd_sc_hs__fa_4 _7637_ (.A(_3450_),
    .B(_3451_),
    .CIN(_3212_),
    .COUT(_3484_),
    .SUM(_3485_));
 sky130_fd_sc_hs__fa_1 _7638_ (.A(_3486_),
    .B(_3487_),
    .CIN(_3488_),
    .COUT(_3489_),
    .SUM(_3490_));
 sky130_fd_sc_hs__fa_1 _7639_ (.A(_3491_),
    .B(_3492_),
    .CIN(_3493_),
    .COUT(_3494_),
    .SUM(_3495_));
 sky130_fd_sc_hs__fa_1 _7640_ (.A(_3496_),
    .B(_3497_),
    .CIN(_3498_),
    .COUT(_3499_),
    .SUM(_3500_));
 sky130_fd_sc_hs__fa_1 _7641_ (.A(_3501_),
    .B(_3502_),
    .CIN(_3503_),
    .COUT(_3504_),
    .SUM(_3505_));
 sky130_fd_sc_hs__fa_1 _7642_ (.A(_3506_),
    .B(_3454_),
    .CIN(_3507_),
    .COUT(_3508_),
    .SUM(_3509_));
 sky130_fd_sc_hs__fa_1 _7643_ (.A(_3510_),
    .B(_3472_),
    .CIN(_3509_),
    .COUT(_3511_),
    .SUM(_3512_));
 sky130_fd_sc_hs__fa_1 _7644_ (.A(_3513_),
    .B(_2778_),
    .CIN(_2779_),
    .COUT(_3514_),
    .SUM(_3515_));
 sky130_fd_sc_hs__fa_1 _7645_ (.A(_3478_),
    .B(_3515_),
    .CIN(_2973_),
    .COUT(_3516_),
    .SUM(_3517_));
 sky130_fd_sc_hs__fa_1 _7646_ (.A(_3480_),
    .B(_3517_),
    .CIN(_3213_),
    .COUT(_3518_),
    .SUM(_3519_));
 sky130_fd_sc_hs__fa_1 _7647_ (.A(_3482_),
    .B(_3519_),
    .CIN(_3485_),
    .COUT(_3520_),
    .SUM(_3521_));
 sky130_fd_sc_hs__fa_1 _7648_ (.A(_3522_),
    .B(_3523_),
    .CIN(_3493_),
    .COUT(_3524_),
    .SUM(_3525_));
 sky130_fd_sc_hs__fa_1 _7649_ (.A(_3526_),
    .B(_3527_),
    .CIN(_3498_),
    .COUT(_3528_),
    .SUM(_3529_));
 sky130_fd_sc_hs__fa_1 _7650_ (.A(_3530_),
    .B(_3531_),
    .CIN(_3532_),
    .COUT(_3533_),
    .SUM(_3534_));
 sky130_fd_sc_hs__fa_1 _7651_ (.A(_3535_),
    .B(_3536_),
    .CIN(_3521_),
    .COUT(_3537_),
    .SUM(_3538_));
 sky130_fd_sc_hs__fa_1 _7652_ (.A(_3539_),
    .B(_3508_),
    .CIN(_3538_),
    .COUT(_3540_),
    .SUM(_3541_));
 sky130_fd_sc_hs__fa_1 _7653_ (.A(_3542_),
    .B(_2778_),
    .CIN(_2779_),
    .COUT(_3543_),
    .SUM(_3544_));
 sky130_fd_sc_hs__fa_1 _7654_ (.A(_3514_),
    .B(_3544_),
    .CIN(_2973_),
    .COUT(_3545_),
    .SUM(_3546_));
 sky130_fd_sc_hs__fa_1 _7655_ (.A(_3516_),
    .B(_3546_),
    .CIN(_3213_),
    .COUT(_3547_),
    .SUM(_3548_));
 sky130_fd_sc_hs__fa_1 _7656_ (.A(_3518_),
    .B(_3548_),
    .CIN(_3485_),
    .COUT(_3549_),
    .SUM(_3550_));
 sky130_fd_sc_hs__fa_2 _7657_ (.A(_3551_),
    .B(_3523_),
    .CIN(_3493_),
    .COUT(_3552_),
    .SUM(_3553_));
 sky130_fd_sc_hs__fa_1 _7658_ (.A(_3524_),
    .B(_3553_),
    .CIN(_3447_),
    .COUT(_3554_),
    .SUM(_3555_));
 sky130_fd_sc_hs__fa_1 _7659_ (.A(_3556_),
    .B(_3557_),
    .CIN(_3532_),
    .COUT(_3558_),
    .SUM(_3559_));
 sky130_fd_sc_hs__fa_1 _7660_ (.A(_3560_),
    .B(_3520_),
    .CIN(_3550_),
    .COUT(_3561_),
    .SUM(_3562_));
 sky130_fd_sc_hs__fa_1 _7661_ (.A(_3563_),
    .B(_3537_),
    .CIN(_3562_),
    .COUT(_3564_),
    .SUM(_3565_));
 sky130_fd_sc_hs__ha_2 _7662_ (.A(_3566_),
    .B(_3567_),
    .COUT(_3568_),
    .SUM(_3569_));
 sky130_fd_sc_hs__ha_4 _7663_ (.A(_3566_),
    .B(net75),
    .COUT(_3570_),
    .SUM(_3571_));
 sky130_fd_sc_hs__ha_1 _7664_ (.A(net74),
    .B(_3567_),
    .COUT(_3572_),
    .SUM(_3573_));
 sky130_fd_sc_hs__ha_4 _7665_ (.A(net74),
    .B(net75),
    .COUT(_3574_),
    .SUM(_3575_));
 sky130_fd_sc_hs__ha_1 _7666_ (.A(_2227_),
    .B(_2228_),
    .COUT(_3576_),
    .SUM(_3577_));
 sky130_fd_sc_hs__ha_4 _7667_ (.A(_3578_),
    .B(_3579_),
    .COUT(_3580_),
    .SUM(_3581_));
 sky130_fd_sc_hs__ha_4 _7668_ (.A(_3582_),
    .B(_3583_),
    .COUT(_3584_),
    .SUM(_3585_));
 sky130_fd_sc_hs__ha_4 _7669_ (.A(_3586_),
    .B(_3587_),
    .COUT(_3588_),
    .SUM(_3589_));
 sky130_fd_sc_hs__ha_4 _7670_ (.A(_3590_),
    .B(_3591_),
    .COUT(_3592_),
    .SUM(_3593_));
 sky130_fd_sc_hs__ha_4 _7671_ (.A(_3594_),
    .B(_3595_),
    .COUT(_3596_),
    .SUM(_3597_));
 sky130_fd_sc_hs__ha_4 _7672_ (.A(_3598_),
    .B(_3599_),
    .COUT(_3600_),
    .SUM(_3601_));
 sky130_fd_sc_hs__ha_4 _7673_ (.A(_3602_),
    .B(_3603_),
    .COUT(_3604_),
    .SUM(_3605_));
 sky130_fd_sc_hs__ha_4 _7674_ (.A(_3606_),
    .B(_3607_),
    .COUT(_3608_),
    .SUM(_3609_));
 sky130_fd_sc_hs__ha_4 _7675_ (.A(_3610_),
    .B(_3611_),
    .COUT(_3612_),
    .SUM(_3613_));
 sky130_fd_sc_hs__ha_2 _7676_ (.A(_3614_),
    .B(_3615_),
    .COUT(_3616_),
    .SUM(_3617_));
 sky130_fd_sc_hs__ha_4 _7677_ (.A(_3618_),
    .B(_3619_),
    .COUT(_3620_),
    .SUM(_3621_));
 sky130_fd_sc_hs__ha_4 _7678_ (.A(_3622_),
    .B(_3623_),
    .COUT(_3624_),
    .SUM(_3625_));
 sky130_fd_sc_hs__ha_4 _7679_ (.A(_3626_),
    .B(_3627_),
    .COUT(_3628_),
    .SUM(_3629_));
 sky130_fd_sc_hs__ha_2 _7680_ (.A(_3630_),
    .B(_3631_),
    .COUT(_3632_),
    .SUM(_3633_));
 sky130_fd_sc_hs__ha_4 _7681_ (.A(_3634_),
    .B(_3635_),
    .COUT(_3636_),
    .SUM(_3637_));
 sky130_fd_sc_hs__ha_1 _7682_ (.A(_3638_),
    .B(_3639_),
    .COUT(_3640_),
    .SUM(_3641_));
 sky130_fd_sc_hs__ha_4 _7683_ (.A(_3642_),
    .B(_3643_),
    .COUT(_3644_),
    .SUM(_3645_));
 sky130_fd_sc_hs__ha_2 _7684_ (.A(_3646_),
    .B(_3647_),
    .COUT(_3648_),
    .SUM(_3649_));
 sky130_fd_sc_hs__ha_2 _7685_ (.A(_3650_),
    .B(_3651_),
    .COUT(_3652_),
    .SUM(_3653_));
 sky130_fd_sc_hs__ha_4 _7686_ (.A(_3654_),
    .B(_3655_),
    .COUT(_3656_),
    .SUM(_3657_));
 sky130_fd_sc_hs__ha_4 _7687_ (.A(_3658_),
    .B(_3659_),
    .COUT(_3660_),
    .SUM(_3661_));
 sky130_fd_sc_hs__ha_2 _7688_ (.A(_3662_),
    .B(_3663_),
    .COUT(_3664_),
    .SUM(_3665_));
 sky130_fd_sc_hs__ha_4 _7689_ (.A(_3666_),
    .B(_3667_),
    .COUT(_3668_),
    .SUM(_3669_));
 sky130_fd_sc_hs__ha_4 _7690_ (.A(_3670_),
    .B(_3671_),
    .COUT(_3672_),
    .SUM(_3673_));
 sky130_fd_sc_hs__ha_4 _7691_ (.A(_3674_),
    .B(_3675_),
    .COUT(_3676_),
    .SUM(_3677_));
 sky130_fd_sc_hs__ha_2 _7692_ (.A(_3678_),
    .B(_3679_),
    .COUT(_3680_),
    .SUM(_3681_));
 sky130_fd_sc_hs__ha_4 _7693_ (.A(_3682_),
    .B(_3683_),
    .COUT(_3684_),
    .SUM(_3685_));
 sky130_fd_sc_hs__ha_2 _7694_ (.A(_3686_),
    .B(_3687_),
    .COUT(_3688_),
    .SUM(_3689_));
 sky130_fd_sc_hs__ha_2 _7695_ (.A(_3690_),
    .B(_3691_),
    .COUT(_3692_),
    .SUM(_3693_));
 sky130_fd_sc_hs__ha_4 _7696_ (.A(_3694_),
    .B(_3695_),
    .COUT(_3696_),
    .SUM(_3697_));
 sky130_fd_sc_hs__ha_4 _7697_ (.A(_3698_),
    .B(_3699_),
    .COUT(_3700_),
    .SUM(_3701_));
 sky130_fd_sc_hs__ha_1 _7698_ (.A(_3702_),
    .B(_3703_),
    .COUT(_3704_),
    .SUM(_3705_));
 sky130_fd_sc_hs__ha_4 _7699_ (.A(_3702_),
    .B(_3703_),
    .COUT(_3706_),
    .SUM(_3707_));
 sky130_fd_sc_hs__ha_1 _7700_ (.A(_3702_),
    .B(\genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .COUT(_3708_),
    .SUM(_3709_));
 sky130_fd_sc_hs__ha_1 _7701_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .B(_3703_),
    .COUT(_3710_),
    .SUM(_3711_));
 sky130_fd_sc_hs__ha_1 _7702_ (.A(\genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .B(\genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .COUT(_3712_),
    .SUM(_3713_));
 sky130_fd_sc_hs__ha_4 _7703_ (.A(_3700_),
    .B(_3714_),
    .COUT(_3715_),
    .SUM(_3716_));
 sky130_fd_sc_hs__ha_4 _7704_ (.A(_3715_),
    .B(_2244_),
    .COUT(_3717_),
    .SUM(_3718_));
 sky130_fd_sc_hs__ha_1 _7705_ (.A(_3719_),
    .B(_3720_),
    .COUT(_2269_),
    .SUM(_3721_));
 sky130_fd_sc_hs__ha_1 _7706_ (.A(_2243_),
    .B(_3722_),
    .COUT(_3723_),
    .SUM(_3724_));
 sky130_fd_sc_hs__ha_1 _7707_ (.A(_3717_),
    .B(_3724_),
    .COUT(_3725_),
    .SUM(_3726_));
 sky130_fd_sc_hs__ha_1 _7708_ (.A(_3723_),
    .B(_2273_),
    .COUT(_3727_),
    .SUM(_3728_));
 sky130_fd_sc_hs__ha_4 _7709_ (.A(_3725_),
    .B(_3728_),
    .COUT(_3729_),
    .SUM(_3730_));
 sky130_fd_sc_hs__ha_1 _7710_ (.A(_3731_),
    .B(_2262_),
    .COUT(_2312_),
    .SUM(_3732_));
 sky130_fd_sc_hs__ha_1 _7711_ (.A(_2272_),
    .B(_3733_),
    .COUT(_3734_),
    .SUM(_3735_));
 sky130_fd_sc_hs__ha_1 _7712_ (.A(_3727_),
    .B(_3735_),
    .COUT(_3736_),
    .SUM(_3737_));
 sky130_fd_sc_hs__ha_4 _7713_ (.A(_3729_),
    .B(_3737_),
    .COUT(_3738_),
    .SUM(_3739_));
 sky130_fd_sc_hs__ha_1 _7714_ (.A(_3740_),
    .B(_3741_),
    .COUT(_2333_),
    .SUM(_3742_));
 sky130_fd_sc_hs__ha_1 _7715_ (.A(_3742_),
    .B(_3743_),
    .COUT(_2342_),
    .SUM(_3744_));
 sky130_fd_sc_hs__ha_1 _7716_ (.A(_3734_),
    .B(_3745_),
    .COUT(_3746_),
    .SUM(_3747_));
 sky130_fd_sc_hs__ha_2 _7717_ (.A(_3736_),
    .B(_3747_),
    .COUT(_2344_),
    .SUM(_3748_));
 sky130_fd_sc_hs__ha_2 _7718_ (.A(_3738_),
    .B(_3748_),
    .COUT(_2343_),
    .SUM(_3749_));
 sky130_fd_sc_hs__ha_1 _7719_ (.A(_3750_),
    .B(_3751_),
    .COUT(_3752_),
    .SUM(_3753_));
 sky130_fd_sc_hs__ha_1 _7720_ (.A(_3746_),
    .B(_3753_),
    .COUT(_3754_),
    .SUM(_2345_));
 sky130_fd_sc_hs__ha_1 _7721_ (.A(_2344_),
    .B(_2345_),
    .COUT(_3755_),
    .SUM(_3756_));
 sky130_fd_sc_hs__ha_1 _7722_ (.A(_3757_),
    .B(_2334_),
    .COUT(_2407_),
    .SUM(_3758_));
 sky130_fd_sc_hs__ha_1 _7723_ (.A(_3759_),
    .B(_3760_),
    .COUT(_3761_),
    .SUM(_3762_));
 sky130_fd_sc_hs__ha_1 _7724_ (.A(_3752_),
    .B(_3762_),
    .COUT(_3763_),
    .SUM(_3764_));
 sky130_fd_sc_hs__ha_4 _7725_ (.A(_3754_),
    .B(_3764_),
    .COUT(_3765_),
    .SUM(_3766_));
 sky130_fd_sc_hs__ha_2 _7726_ (.A(_3767_),
    .B(_3768_),
    .COUT(_3769_),
    .SUM(_3770_));
 sky130_fd_sc_hs__ha_1 _7727_ (.A(_3770_),
    .B(_2368_),
    .COUT(_3771_),
    .SUM(_3772_));
 sky130_fd_sc_hs__ha_2 _7728_ (.A(_3761_),
    .B(_3773_),
    .COUT(_3774_),
    .SUM(_3775_));
 sky130_fd_sc_hs__ha_4 _7729_ (.A(_3763_),
    .B(_3775_),
    .COUT(_3776_),
    .SUM(_3777_));
 sky130_fd_sc_hs__ha_1 _7730_ (.A(_3769_),
    .B(_2439_),
    .COUT(_2481_),
    .SUM(_3778_));
 sky130_fd_sc_hs__ha_1 _7731_ (.A(_3778_),
    .B(_2396_),
    .COUT(_3779_),
    .SUM(_3780_));
 sky130_fd_sc_hs__ha_1 _7732_ (.A(_3781_),
    .B(_3782_),
    .COUT(_3783_),
    .SUM(_3784_));
 sky130_fd_sc_hs__ha_4 _7733_ (.A(_3774_),
    .B(_3784_),
    .COUT(_3785_),
    .SUM(_3786_));
 sky130_fd_sc_hs__ha_1 _7734_ (.A(_3787_),
    .B(_3788_),
    .COUT(_3789_),
    .SUM(_3790_));
 sky130_fd_sc_hs__ha_2 _7735_ (.A(_3783_),
    .B(_3790_),
    .COUT(_3791_),
    .SUM(_3792_));
 sky130_fd_sc_hs__ha_1 _7736_ (.A(_3793_),
    .B(_3794_),
    .COUT(_3795_),
    .SUM(_3796_));
 sky130_fd_sc_hs__ha_1 _7737_ (.A(_3797_),
    .B(_2536_),
    .COUT(_3798_),
    .SUM(_3799_));
 sky130_fd_sc_hs__ha_2 _7738_ (.A(_3789_),
    .B(_3799_),
    .COUT(_3800_),
    .SUM(_3801_));
 sky130_fd_sc_hs__ha_1 _7739_ (.A(_3795_),
    .B(_3802_),
    .COUT(_2649_),
    .SUM(_2587_));
 sky130_fd_sc_hs__ha_1 _7740_ (.A(_2535_),
    .B(_2591_),
    .COUT(_3803_),
    .SUM(_3804_));
 sky130_fd_sc_hs__ha_4 _7741_ (.A(_3798_),
    .B(_3804_),
    .COUT(_3805_),
    .SUM(_3806_));
 sky130_fd_sc_hs__ha_1 _7742_ (.A(_3807_),
    .B(_2572_),
    .COUT(_3808_),
    .SUM(_3809_));
 sky130_fd_sc_hs__ha_1 _7743_ (.A(_3809_),
    .B(_2582_),
    .COUT(_2702_),
    .SUM(_3810_));
 sky130_fd_sc_hs__ha_4 _7744_ (.A(_3803_),
    .B(_3811_),
    .COUT(_3812_),
    .SUM(_3813_));
 sky130_fd_sc_hs__ha_1 _7745_ (.A(_3814_),
    .B(_3815_),
    .COUT(_2754_),
    .SUM(_3816_));
 sky130_fd_sc_hs__ha_1 _7746_ (.A(_3816_),
    .B(_2627_),
    .COUT(_3817_),
    .SUM(_3818_));
 sky130_fd_sc_hs__ha_1 _7747_ (.A(_3808_),
    .B(_3818_),
    .COUT(_2762_),
    .SUM(_3819_));
 sky130_fd_sc_hs__ha_1 _7748_ (.A(_3819_),
    .B(_2637_),
    .COUT(_2773_),
    .SUM(_3820_));
 sky130_fd_sc_hs__ha_4 _7749_ (.A(_3821_),
    .B(_3822_),
    .COUT(_3823_),
    .SUM(_3824_));
 sky130_fd_sc_hs__ha_4 _7750_ (.A(_3825_),
    .B(_3826_),
    .COUT(_3827_),
    .SUM(_3828_));
 sky130_fd_sc_hs__ha_1 _7751_ (.A(_2755_),
    .B(_3829_),
    .COUT(_2893_),
    .SUM(_3830_));
 sky130_fd_sc_hs__ha_2 _7752_ (.A(_3831_),
    .B(_3832_),
    .COUT(_3833_),
    .SUM(_3834_));
 sky130_fd_sc_hs__ha_1 _7753_ (.A(_3835_),
    .B(_3836_),
    .COUT(_2956_),
    .SUM(_2894_));
 sky130_fd_sc_hs__ha_4 _7754_ (.A(_3837_),
    .B(_3838_),
    .COUT(_3839_),
    .SUM(_3840_));
 sky130_fd_sc_hs__ha_1 _7755_ (.A(_3841_),
    .B(_3842_),
    .COUT(_3019_),
    .SUM(_2957_));
 sky130_fd_sc_hs__ha_2 _7756_ (.A(_3843_),
    .B(_3844_),
    .COUT(_3845_),
    .SUM(_3846_));
 sky130_fd_sc_hs__ha_1 _7757_ (.A(_3847_),
    .B(_3848_),
    .COUT(_3078_),
    .SUM(_3020_));
 sky130_fd_sc_hs__ha_4 _7758_ (.A(_3849_),
    .B(_3850_),
    .COUT(_3851_),
    .SUM(_3852_));
 sky130_fd_sc_hs__ha_1 _7759_ (.A(_3853_),
    .B(_3854_),
    .COUT(_3135_),
    .SUM(_3079_));
 sky130_fd_sc_hs__ha_4 _7760_ (.A(_3855_),
    .B(_3856_),
    .COUT(_3857_),
    .SUM(_3858_));
 sky130_fd_sc_hs__ha_1 _7761_ (.A(_3859_),
    .B(_3860_),
    .COUT(_3193_),
    .SUM(_3136_));
 sky130_fd_sc_hs__ha_2 _7762_ (.A(_3861_),
    .B(_3862_),
    .COUT(_3863_),
    .SUM(_3864_));
 sky130_fd_sc_hs__ha_1 _7763_ (.A(_3865_),
    .B(_3866_),
    .COUT(_3247_),
    .SUM(_3194_));
 sky130_fd_sc_hs__ha_2 _7764_ (.A(_3867_),
    .B(_3868_),
    .COUT(_3869_),
    .SUM(_3870_));
 sky130_fd_sc_hs__ha_1 _7765_ (.A(_3871_),
    .B(_3872_),
    .COUT(_3297_),
    .SUM(_3248_));
 sky130_fd_sc_hs__ha_2 _7766_ (.A(_3873_),
    .B(_3874_),
    .COUT(_3875_),
    .SUM(_3876_));
 sky130_fd_sc_hs__ha_1 _7767_ (.A(_3877_),
    .B(_3878_),
    .COUT(_3346_),
    .SUM(_3298_));
 sky130_fd_sc_hs__ha_2 _7768_ (.A(_3879_),
    .B(_3880_),
    .COUT(_3881_),
    .SUM(_3882_));
 sky130_fd_sc_hs__ha_1 _7769_ (.A(_3883_),
    .B(_3884_),
    .COUT(_3389_),
    .SUM(_3347_));
 sky130_fd_sc_hs__ha_2 _7770_ (.A(_3885_),
    .B(_3886_),
    .COUT(_3887_),
    .SUM(_3888_));
 sky130_fd_sc_hs__ha_1 _7771_ (.A(_3889_),
    .B(_3890_),
    .COUT(_3428_),
    .SUM(_3390_));
 sky130_fd_sc_hs__ha_2 _7772_ (.A(_3891_),
    .B(_3892_),
    .COUT(_3893_),
    .SUM(_3894_));
 sky130_fd_sc_hs__ha_1 _7773_ (.A(_3895_),
    .B(_3896_),
    .COUT(_3466_),
    .SUM(_3429_));
 sky130_fd_sc_hs__ha_4 _7774_ (.A(_3897_),
    .B(_3898_),
    .COUT(_3899_),
    .SUM(_3900_));
 sky130_fd_sc_hs__ha_1 _7775_ (.A(_3901_),
    .B(_3902_),
    .COUT(_3501_),
    .SUM(_3467_));
 sky130_fd_sc_hs__ha_2 _7776_ (.A(_3903_),
    .B(_3904_),
    .COUT(_3905_),
    .SUM(_3906_));
 sky130_fd_sc_hs__ha_1 _7777_ (.A(_3907_),
    .B(_3908_),
    .COUT(_3530_),
    .SUM(_3502_));
 sky130_fd_sc_hs__ha_2 _7778_ (.A(_3909_),
    .B(_3910_),
    .COUT(_3911_),
    .SUM(_3912_));
 sky130_fd_sc_hs__ha_1 _7779_ (.A(_3913_),
    .B(_3914_),
    .COUT(_3556_),
    .SUM(_3531_));
 sky130_fd_sc_hs__ha_4 _7780_ (.A(_3915_),
    .B(_3916_),
    .COUT(_3917_),
    .SUM(_3918_));
 sky130_fd_sc_hs__ha_1 _7781_ (.A(_3553_),
    .B(_3447_),
    .COUT(_3919_),
    .SUM(_3920_));
 sky130_fd_sc_hs__ha_1 _7782_ (.A(_3921_),
    .B(_3555_),
    .COUT(_3922_),
    .SUM(_3557_));
 sky130_fd_sc_hs__ha_4 _7783_ (.A(_3923_),
    .B(_3924_),
    .COUT(_3925_),
    .SUM(_3926_));
 sky130_fd_sc_hs__ha_4 _7784_ (.A(_3927_),
    .B(_3928_),
    .COUT(_3929_),
    .SUM(_3930_));
 sky130_fd_sc_hs__ha_1 _7785_ (.A(net34),
    .B(net66),
    .COUT(_3931_),
    .SUM(_3932_));
 sky130_fd_sc_hs__ha_2 _7786_ (.A(_3933_),
    .B(_3934_),
    .COUT(_3935_),
    .SUM(_3936_));
 sky130_fd_sc_hs__ha_1 _7787_ (.A(_3937_),
    .B(_3933_),
    .COUT(_3938_),
    .SUM(_3939_));
 sky130_fd_sc_hs__ha_1 _7788_ (.A(net2),
    .B(net42),
    .COUT(_3940_),
    .SUM(_3941_));
 sky130_fd_sc_hs__ha_1 _7789_ (.A(_3942_),
    .B(_3934_),
    .COUT(_3943_),
    .SUM(_3944_));
 sky130_fd_sc_hs__ha_1 _7790_ (.A(net21),
    .B(net53),
    .COUT(_3945_),
    .SUM(_3946_));
 sky130_fd_sc_hs__ha_1 _7791_ (.A(_3947_),
    .B(_3948_),
    .COUT(_3949_),
    .SUM(_3950_));
 sky130_fd_sc_hs__ha_1 _7792_ (.A(net32),
    .B(net64),
    .COUT(_3951_),
    .SUM(_3952_));
 sky130_fd_sc_hs__ha_1 _7793_ (.A(_3953_),
    .B(_3954_),
    .COUT(_3955_),
    .SUM(_3956_));
 sky130_fd_sc_hs__ha_1 _7794_ (.A(net35),
    .B(net67),
    .COUT(_3957_),
    .SUM(_3958_));
 sky130_fd_sc_hs__ha_1 _7795_ (.A(_3959_),
    .B(_3960_),
    .COUT(_3961_),
    .SUM(_3962_));
 sky130_fd_sc_hs__ha_1 _7796_ (.A(net36),
    .B(net68),
    .COUT(_3963_),
    .SUM(_3964_));
 sky130_fd_sc_hs__ha_1 _7797_ (.A(_3965_),
    .B(_3966_),
    .COUT(_3967_),
    .SUM(_3968_));
 sky130_fd_sc_hs__ha_1 _7798_ (.A(net37),
    .B(net69),
    .COUT(_3969_),
    .SUM(_3970_));
 sky130_fd_sc_hs__ha_1 _7799_ (.A(_3971_),
    .B(_3972_),
    .COUT(_3973_),
    .SUM(_3974_));
 sky130_fd_sc_hs__ha_1 _7800_ (.A(net38),
    .B(net70),
    .COUT(_3975_),
    .SUM(_3976_));
 sky130_fd_sc_hs__ha_1 _7801_ (.A(_3977_),
    .B(_3978_),
    .COUT(_3979_),
    .SUM(_3980_));
 sky130_fd_sc_hs__ha_1 _7802_ (.A(net39),
    .B(net71),
    .COUT(_3981_),
    .SUM(_3982_));
 sky130_fd_sc_hs__ha_1 _7803_ (.A(_3983_),
    .B(_3984_),
    .COUT(_3985_),
    .SUM(_3986_));
 sky130_fd_sc_hs__ha_1 _7804_ (.A(net40),
    .B(net72),
    .COUT(_3987_),
    .SUM(_3988_));
 sky130_fd_sc_hs__ha_1 _7805_ (.A(_3989_),
    .B(_3990_),
    .COUT(_3991_),
    .SUM(_3992_));
 sky130_fd_sc_hs__ha_1 _7806_ (.A(net41),
    .B(net73),
    .COUT(_3993_),
    .SUM(_3994_));
 sky130_fd_sc_hs__ha_1 _7807_ (.A(_3995_),
    .B(_3996_),
    .COUT(_3997_),
    .SUM(_3998_));
 sky130_fd_sc_hs__ha_1 _7808_ (.A(net3),
    .B(net43),
    .COUT(_3999_),
    .SUM(_4000_));
 sky130_fd_sc_hs__ha_1 _7809_ (.A(_4001_),
    .B(_4002_),
    .COUT(_4003_),
    .SUM(_4004_));
 sky130_fd_sc_hs__ha_1 _7810_ (.A(net4),
    .B(net44),
    .COUT(_4005_),
    .SUM(_4006_));
 sky130_fd_sc_hs__ha_1 _7811_ (.A(_4007_),
    .B(_4008_),
    .COUT(_4009_),
    .SUM(_4010_));
 sky130_fd_sc_hs__ha_1 _7812_ (.A(net5),
    .B(net45),
    .COUT(_4011_),
    .SUM(_4012_));
 sky130_fd_sc_hs__ha_1 _7813_ (.A(_4013_),
    .B(_4014_),
    .COUT(_4015_),
    .SUM(_4016_));
 sky130_fd_sc_hs__ha_1 _7814_ (.A(net6),
    .B(net46),
    .COUT(_4017_),
    .SUM(_4018_));
 sky130_fd_sc_hs__ha_1 _7815_ (.A(_4019_),
    .B(_4020_),
    .COUT(_4021_),
    .SUM(_4022_));
 sky130_fd_sc_hs__ha_1 _7816_ (.A(net7),
    .B(net47),
    .COUT(_4023_),
    .SUM(_4024_));
 sky130_fd_sc_hs__ha_1 _7817_ (.A(_4025_),
    .B(_4026_),
    .COUT(_4027_),
    .SUM(_4028_));
 sky130_fd_sc_hs__ha_1 _7818_ (.A(net8),
    .B(net48),
    .COUT(_4029_),
    .SUM(_4030_));
 sky130_fd_sc_hs__ha_1 _7819_ (.A(_4031_),
    .B(_4032_),
    .COUT(_4033_),
    .SUM(_4034_));
 sky130_fd_sc_hs__ha_1 _7820_ (.A(net17),
    .B(net49),
    .COUT(_4035_),
    .SUM(_4036_));
 sky130_fd_sc_hs__ha_1 _7821_ (.A(_4037_),
    .B(_4038_),
    .COUT(_4039_),
    .SUM(_4040_));
 sky130_fd_sc_hs__ha_1 _7822_ (.A(net18),
    .B(net50),
    .COUT(_4041_),
    .SUM(_4042_));
 sky130_fd_sc_hs__ha_1 _7823_ (.A(_4043_),
    .B(_4044_),
    .COUT(_4045_),
    .SUM(_4046_));
 sky130_fd_sc_hs__ha_1 _7824_ (.A(net19),
    .B(net51),
    .COUT(_4047_),
    .SUM(_4048_));
 sky130_fd_sc_hs__ha_1 _7825_ (.A(_4049_),
    .B(_4050_),
    .COUT(_4051_),
    .SUM(_4052_));
 sky130_fd_sc_hs__ha_1 _7826_ (.A(net20),
    .B(net52),
    .COUT(_4053_),
    .SUM(_4054_));
 sky130_fd_sc_hs__ha_1 _7827_ (.A(_4055_),
    .B(_4056_),
    .COUT(_4057_),
    .SUM(_4058_));
 sky130_fd_sc_hs__ha_1 _7828_ (.A(net22),
    .B(net54),
    .COUT(_4059_),
    .SUM(_4060_));
 sky130_fd_sc_hs__ha_1 _7829_ (.A(_4061_),
    .B(_4062_),
    .COUT(_4063_),
    .SUM(_4064_));
 sky130_fd_sc_hs__ha_1 _7830_ (.A(net23),
    .B(net55),
    .COUT(_4065_),
    .SUM(_4066_));
 sky130_fd_sc_hs__ha_1 _7831_ (.A(_4067_),
    .B(_4068_),
    .COUT(_4069_),
    .SUM(_4070_));
 sky130_fd_sc_hs__ha_1 _7832_ (.A(net24),
    .B(net56),
    .COUT(_4071_),
    .SUM(_4072_));
 sky130_fd_sc_hs__ha_1 _7833_ (.A(_4073_),
    .B(_4074_),
    .COUT(_4075_),
    .SUM(_4076_));
 sky130_fd_sc_hs__ha_1 _7834_ (.A(net25),
    .B(net57),
    .COUT(_4077_),
    .SUM(_4078_));
 sky130_fd_sc_hs__ha_1 _7835_ (.A(_4079_),
    .B(_4080_),
    .COUT(_4081_),
    .SUM(_4082_));
 sky130_fd_sc_hs__ha_1 _7836_ (.A(net26),
    .B(net58),
    .COUT(_4083_),
    .SUM(_4084_));
 sky130_fd_sc_hs__ha_1 _7837_ (.A(_4085_),
    .B(_4086_),
    .COUT(_4087_),
    .SUM(_4088_));
 sky130_fd_sc_hs__ha_1 _7838_ (.A(net27),
    .B(net59),
    .COUT(_4089_),
    .SUM(_4090_));
 sky130_fd_sc_hs__ha_1 _7839_ (.A(_4091_),
    .B(_4092_),
    .COUT(_4093_),
    .SUM(_4094_));
 sky130_fd_sc_hs__ha_1 _7840_ (.A(net28),
    .B(net60),
    .COUT(_4095_),
    .SUM(_4096_));
 sky130_fd_sc_hs__ha_1 _7841_ (.A(_4097_),
    .B(_4098_),
    .COUT(_4099_),
    .SUM(_4100_));
 sky130_fd_sc_hs__ha_1 _7842_ (.A(net29),
    .B(net61),
    .COUT(_4101_),
    .SUM(_4102_));
 sky130_fd_sc_hs__ha_1 _7843_ (.A(_4103_),
    .B(_4104_),
    .COUT(_4105_),
    .SUM(_4106_));
 sky130_fd_sc_hs__ha_1 _7844_ (.A(net30),
    .B(net62),
    .COUT(_4107_),
    .SUM(_4108_));
 sky130_fd_sc_hs__ha_1 _7845_ (.A(_4109_),
    .B(_4110_),
    .COUT(_4111_),
    .SUM(_4112_));
 sky130_fd_sc_hs__ha_1 _7846_ (.A(net31),
    .B(net63),
    .COUT(_4113_),
    .SUM(_4114_));
 sky130_fd_sc_hs__ha_1 _7847_ (.A(_4115_),
    .B(_4116_),
    .COUT(_4117_),
    .SUM(_4118_));
 sky130_fd_sc_hs__ha_1 _7848_ (.A(net33),
    .B(net65),
    .COUT(_4119_),
    .SUM(_4120_));
 sky130_fd_sc_hs__dfrtp_1 _7849_ (.D(_0006_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[2] ),
    .RESET_B(net357),
    .CLK(clknet_3_0_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 _7850_ (.D(_0007_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[1] ),
    .RESET_B(net357),
    .CLK(clknet_3_0_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 _7851_ (.D(_0008_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.md_state_q[5] ),
    .RESET_B(net360),
    .CLK(clknet_3_1_0_clk_i));
 sky130_fd_sc_hs__dfrtp_2 _7852_ (.D(_0009_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.md_state_q[2] ),
    .RESET_B(net359),
    .CLK(clknet_3_1_0_clk_i));
 sky130_fd_sc_hs__dfstp_1 _7853_ (.D(_0010_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.md_state_q[0] ),
    .SET_B(net360),
    .CLK(clknet_3_1_0_clk_i));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_0_clk_i (.A(clk_i),
    .X(clknet_0_clk_i));
 sky130_fd_sc_hs__buf_8 _7855_ (.A(net191),
    .X(net224));
 sky130_fd_sc_hs__clkbuf_4 _7856_ (.A(net202),
    .X(net235));
 sky130_fd_sc_hs__buf_8 _7857_ (.A(net213),
    .X(net246));
 sky130_fd_sc_hs__buf_4 _7858_ (.A(net216),
    .X(net249));
 sky130_fd_sc_hs__buf_8 _7859_ (.A(net217),
    .X(net250));
 sky130_fd_sc_hs__clkbuf_4 _7860_ (.A(net218),
    .X(net251));
 sky130_fd_sc_hs__clkbuf_8 _7861_ (.A(net219),
    .X(net252));
 sky130_fd_sc_hs__buf_8 _7862_ (.A(net220),
    .X(net253));
 sky130_fd_sc_hs__buf_8 _7863_ (.A(net221),
    .X(net254));
 sky130_fd_sc_hs__clkbuf_4 _7864_ (.A(net222),
    .X(net255));
 sky130_fd_sc_hs__buf_4 _7865_ (.A(net192),
    .X(net225));
 sky130_fd_sc_hs__buf_8 _7866_ (.A(net193),
    .X(net226));
 sky130_fd_sc_hs__buf_2 _7867_ (.A(net194),
    .X(net227));
 sky130_fd_sc_hs__buf_8 _7868_ (.A(net195),
    .X(net228));
 sky130_fd_sc_hs__clkbuf_8 _7869_ (.A(net16),
    .X(net229));
 sky130_fd_sc_hs__buf_4 _7870_ (.A(net197),
    .X(net230));
 sky130_fd_sc_hs__clkbuf_8 _7871_ (.A(net198),
    .X(net231));
 sky130_fd_sc_hs__clkbuf_8 _7872_ (.A(net199),
    .X(net232));
 sky130_fd_sc_hs__clkbuf_8 _7873_ (.A(net200),
    .X(net233));
 sky130_fd_sc_hs__buf_4 _7874_ (.A(net201),
    .X(net234));
 sky130_fd_sc_hs__buf_8 _7875_ (.A(net203),
    .X(net236));
 sky130_fd_sc_hs__buf_4 _7876_ (.A(net204),
    .X(net237));
 sky130_fd_sc_hs__buf_8 _7877_ (.A(net205),
    .X(net238));
 sky130_fd_sc_hs__buf_8 _7878_ (.A(net206),
    .X(net239));
 sky130_fd_sc_hs__buf_4 _7879_ (.A(net207),
    .X(net240));
 sky130_fd_sc_hs__buf_8 _7880_ (.A(net208),
    .X(net241));
 sky130_fd_sc_hs__buf_8 _7881_ (.A(net209),
    .X(net242));
 sky130_fd_sc_hs__clkbuf_8 _7882_ (.A(net210),
    .X(net243));
 sky130_fd_sc_hs__buf_4 _7883_ (.A(net211),
    .X(net244));
 sky130_fd_sc_hs__buf_4 _7884_ (.A(net212),
    .X(net245));
 sky130_fd_sc_hs__clkbuf_8 _7885_ (.A(net214),
    .X(net247));
 sky130_fd_sc_hs__buf_8 _7886_ (.A(net215),
    .X(net248));
 sky130_fd_sc_hs__buf_4 _7887_ (.A(net363),
    .X(imd_val_d_o[32]));
 sky130_fd_sc_hs__buf_4 _7888_ (.A(net364),
    .X(imd_val_d_o[33]));
 sky130_fd_sc_hs__dfrtp_2 \genblk3.gen_multdiv_fast.multdiv_i.div_by_zero_q$_DFFE_PN0P_  (.D(_0011_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.div_by_zero_q ),
    .RESET_B(net360),
    .CLK(clknet_3_1_0_clk_i));
 sky130_fd_sc_hs__dfrtp_2 \genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0]$_DFFE_PN0P_  (.D(_0012_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[0] ),
    .RESET_B(net360),
    .CLK(clknet_3_3_0_clk_i));
 sky130_fd_sc_hs__dfrtp_2 \genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1]$_DFFE_PN0P_  (.D(_0013_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[1] ),
    .RESET_B(net360),
    .CLK(clknet_3_6_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[2]$_DFFE_PN0P_  (.D(_0014_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[2] ),
    .RESET_B(net360),
    .CLK(clknet_3_3_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[3]$_DFFE_PN0P_  (.D(_0015_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[3] ),
    .RESET_B(net360),
    .CLK(clknet_3_6_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[4]$_DFFE_PN0P_  (.D(_0016_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.div_counter_q[4] ),
    .RESET_B(net360),
    .CLK(clknet_3_3_0_clk_i));
 sky130_fd_sc_hs__dfstp_1 \genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0]$_DFF_PN1_  (.D(_0000_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[0] ),
    .SET_B(net357),
    .CLK(clknet_3_0_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3]$_DFF_PN0_  (.D(_0001_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.gen_mult_fast.mult_state_q[3] ),
    .RESET_B(net357),
    .CLK(clknet_3_0_0_clk_i));
 sky130_fd_sc_hs__dfrtp_2 \genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1]$_DFF_PN0_  (.D(_0002_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.md_state_q[1] ),
    .RESET_B(net360),
    .CLK(clknet_3_1_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.md_state_q[3]$_DFF_PN0_  (.D(_0003_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.div_valid ),
    .RESET_B(net360),
    .CLK(clknet_3_1_0_clk_i));
 sky130_fd_sc_hs__dfrtp_4 \genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4]$_DFF_PN0_  (.D(_0004_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.md_state_q[4] ),
    .RESET_B(net360),
    .CLK(clknet_3_1_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.md_state_q[6]$_DFF_PN0_  (.D(_0005_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.md_state_q[6] ),
    .RESET_B(net360),
    .CLK(clknet_3_1_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[0]$_DFFE_PN0P_  (.D(_0017_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[0] ),
    .RESET_B(net358),
    .CLK(clknet_3_2_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[10]$_DFFE_PN0P_  (.D(_0018_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[10] ),
    .RESET_B(net359),
    .CLK(clknet_3_1_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[11]$_DFFE_PN0P_  (.D(_0019_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[11] ),
    .RESET_B(net359),
    .CLK(clknet_3_3_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[12]$_DFFE_PN0P_  (.D(_0020_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[12] ),
    .RESET_B(net358),
    .CLK(clknet_3_2_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[13]$_DFFE_PN0P_  (.D(_0021_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[13] ),
    .RESET_B(net359),
    .CLK(clknet_3_3_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[14]$_DFFE_PN0P_  (.D(_0022_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[14] ),
    .RESET_B(net359),
    .CLK(clknet_3_3_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[15]$_DFFE_PN0P_  (.D(_0023_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[15] ),
    .RESET_B(net358),
    .CLK(clknet_3_2_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[16]$_DFFE_PN0P_  (.D(_0024_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[16] ),
    .RESET_B(net357),
    .CLK(clknet_3_2_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[17]$_DFFE_PN0P_  (.D(_0025_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[17] ),
    .RESET_B(net357),
    .CLK(clknet_3_2_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[18]$_DFFE_PN0P_  (.D(_0026_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[18] ),
    .RESET_B(net357),
    .CLK(clknet_3_2_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[19]$_DFFE_PN0P_  (.D(_0027_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[19] ),
    .RESET_B(net357),
    .CLK(clknet_3_2_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[1]$_DFFE_PN0P_  (.D(_0028_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[1] ),
    .RESET_B(net358),
    .CLK(clknet_3_0_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[20]$_DFFE_PN0P_  (.D(_0029_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[20] ),
    .RESET_B(net358),
    .CLK(clknet_3_0_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[21]$_DFFE_PN0P_  (.D(_0030_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[21] ),
    .RESET_B(net357),
    .CLK(clknet_3_0_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[22]$_DFFE_PN0P_  (.D(_0031_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[22] ),
    .RESET_B(net357),
    .CLK(clknet_3_0_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[23]$_DFFE_PN0P_  (.D(_0032_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[23] ),
    .RESET_B(net357),
    .CLK(clknet_3_0_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[24]$_DFFE_PN0P_  (.D(_0033_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[24] ),
    .RESET_B(net357),
    .CLK(clknet_3_2_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[25]$_DFFE_PN0P_  (.D(_0034_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[25] ),
    .RESET_B(net357),
    .CLK(clknet_3_2_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[26]$_DFFE_PN0P_  (.D(_0035_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[26] ),
    .RESET_B(net357),
    .CLK(clknet_3_2_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[27]$_DFFE_PN0P_  (.D(_0036_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[27] ),
    .RESET_B(net358),
    .CLK(clknet_3_0_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[28]$_DFFE_PN0P_  (.D(_0037_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[28] ),
    .RESET_B(net358),
    .CLK(clknet_3_0_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[29]$_DFFE_PN0P_  (.D(_0038_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[29] ),
    .RESET_B(net358),
    .CLK(clknet_3_0_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[2]$_DFFE_PN0P_  (.D(_0039_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[2] ),
    .RESET_B(net358),
    .CLK(clknet_3_2_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[30]$_DFFE_PN0P_  (.D(_0040_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[30] ),
    .RESET_B(net358),
    .CLK(clknet_3_0_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[31]$_DFFE_PN0P_  (.D(_0041_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[31] ),
    .RESET_B(net358),
    .CLK(clknet_3_0_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[3]$_DFFE_PN0P_  (.D(_0042_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[3] ),
    .RESET_B(net358),
    .CLK(clknet_3_2_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[4]$_DFFE_PN0P_  (.D(_0043_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[4] ),
    .RESET_B(net359),
    .CLK(clknet_3_1_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[5]$_DFFE_PN0P_  (.D(_0044_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[5] ),
    .RESET_B(net359),
    .CLK(clknet_3_3_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[6]$_DFFE_PN0P_  (.D(_0045_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[6] ),
    .RESET_B(net359),
    .CLK(clknet_3_3_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[7]$_DFFE_PN0P_  (.D(_0046_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[7] ),
    .RESET_B(net359),
    .CLK(clknet_3_3_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[8]$_DFFE_PN0P_  (.D(_0047_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[8] ),
    .RESET_B(net359),
    .CLK(clknet_3_1_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[9]$_DFFE_PN0P_  (.D(_0048_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_numerator_q[9] ),
    .RESET_B(net359),
    .CLK(clknet_3_1_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[0]$_DFFE_PN0P_  (.D(_0049_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[0] ),
    .RESET_B(net361),
    .CLK(clknet_3_7_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[10]$_DFFE_PN0P_  (.D(_0050_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[10] ),
    .RESET_B(net190),
    .CLK(clknet_3_5_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[11]$_DFFE_PN0P_  (.D(_0051_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[11] ),
    .RESET_B(net190),
    .CLK(clknet_3_5_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[12]$_DFFE_PN0P_  (.D(_0052_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[12] ),
    .RESET_B(net362),
    .CLK(clknet_3_5_0_clk_i));
 sky130_fd_sc_hs__dfrtp_2 \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[13]$_DFFE_PN0P_  (.D(_0053_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[13] ),
    .RESET_B(net362),
    .CLK(clknet_3_5_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[14]$_DFFE_PN0P_  (.D(_0054_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[14] ),
    .RESET_B(net190),
    .CLK(clknet_3_5_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[15]$_DFFE_PN0P_  (.D(_0055_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[15] ),
    .RESET_B(net190),
    .CLK(clknet_3_5_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[16]$_DFFE_PN0P_  (.D(_0056_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[16] ),
    .RESET_B(net361),
    .CLK(clknet_3_4_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[17]$_DFFE_PN0P_  (.D(_0057_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[17] ),
    .RESET_B(net362),
    .CLK(clknet_3_5_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[18]$_DFFE_PN0P_  (.D(_0058_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[18] ),
    .RESET_B(net362),
    .CLK(clknet_3_7_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[19]$_DFFE_PN0P_  (.D(_0059_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[19] ),
    .RESET_B(net362),
    .CLK(clknet_3_7_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[1]$_DFFE_PN0P_  (.D(_0060_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[1] ),
    .RESET_B(net361),
    .CLK(clknet_3_4_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[20]$_DFFE_PN0P_  (.D(_0061_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[20] ),
    .RESET_B(net361),
    .CLK(clknet_3_7_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[21]$_DFFE_PN0P_  (.D(_0062_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[21] ),
    .RESET_B(net362),
    .CLK(clknet_3_7_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[22]$_DFFE_PN0P_  (.D(_0063_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[22] ),
    .RESET_B(net362),
    .CLK(clknet_3_7_0_clk_i));
 sky130_fd_sc_hs__dfrtp_2 \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[23]$_DFFE_PN0P_  (.D(_0064_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[23] ),
    .RESET_B(net361),
    .CLK(clknet_3_7_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[24]$_DFFE_PN0P_  (.D(_0065_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[24] ),
    .RESET_B(net362),
    .CLK(clknet_3_4_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[25]$_DFFE_PN0P_  (.D(_0066_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[25] ),
    .RESET_B(net362),
    .CLK(clknet_3_4_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[26]$_DFFE_PN0P_  (.D(_0067_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[26] ),
    .RESET_B(net361),
    .CLK(clknet_3_4_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[27]$_DFFE_PN0P_  (.D(_0068_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[27] ),
    .RESET_B(net361),
    .CLK(clknet_3_4_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[28]$_DFFE_PN0P_  (.D(_0069_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[28] ),
    .RESET_B(net361),
    .CLK(clknet_3_6_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[29]$_DFFE_PN0P_  (.D(_0070_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[29] ),
    .RESET_B(net361),
    .CLK(clknet_3_6_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[2]$_DFFE_PN0P_  (.D(_0071_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[2] ),
    .RESET_B(net361),
    .CLK(clknet_3_6_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[30]$_DFFE_PN0P_  (.D(_0072_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[30] ),
    .RESET_B(net361),
    .CLK(clknet_3_6_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[31]$_DFFE_PN0P_  (.D(_0073_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[31] ),
    .RESET_B(net361),
    .CLK(clknet_3_6_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[3]$_DFFE_PN0P_  (.D(_0074_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[3] ),
    .RESET_B(net361),
    .CLK(clknet_3_6_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[4]$_DFFE_PN0P_  (.D(_0075_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[4] ),
    .RESET_B(net361),
    .CLK(clknet_3_7_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[5]$_DFFE_PN0P_  (.D(_0076_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[5] ),
    .RESET_B(net362),
    .CLK(clknet_3_5_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[6]$_DFFE_PN0P_  (.D(_0077_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[6] ),
    .RESET_B(net362),
    .CLK(clknet_3_7_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[7]$_DFFE_PN0P_  (.D(_0078_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[7] ),
    .RESET_B(net190),
    .CLK(clknet_3_5_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[8]$_DFFE_PN0P_  (.D(_0079_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[8] ),
    .RESET_B(net360),
    .CLK(clknet_3_4_0_clk_i));
 sky130_fd_sc_hs__dfrtp_1 \genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[9]$_DFFE_PN0P_  (.D(_0080_),
    .Q(\genblk3.gen_multdiv_fast.multdiv_i.op_quotient_q[9] ),
    .RESET_B(net362),
    .CLK(clknet_3_5_0_clk_i));
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_7 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_8 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_9 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_10 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_11 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_12 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_13 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_14 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_15 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_16 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_17 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_18 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_19 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_20 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_21 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_22 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_23 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_24 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_25 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_26 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_27 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_28 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_29 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_30 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_31 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_32 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_33 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_34 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_35 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_36 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_37 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_38 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_39 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_40 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_41 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_42 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_43 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_44 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_45 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_46 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_47 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_48 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_49 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_50 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_51 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_52 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_53 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_54 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_55 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_56 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_57 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_58 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_59 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_60 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_61 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_62 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_63 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_64 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_65 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_66 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_67 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_68 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_69 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_70 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_71 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_72 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_73 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_74 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_75 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_76 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_77 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_78 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_79 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_80 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_81 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_82 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_83 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_84 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_85 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_86 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_87 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_88 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_89 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_90 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_91 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_92 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_93 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_94 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_95 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_96 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_97 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_98 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_99 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_100 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_101 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_102 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_103 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_104 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_105 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_106 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_107 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_108 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_109 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_110 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_111 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_112 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_113 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_114 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_115 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_116 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_117 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_118 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_119 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_120 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_121 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_122 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_123 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_124 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_125 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_126 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_127 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_128 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_129 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_130 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_131 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_132 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_133 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_134 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_135 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_136 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_137 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_138 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_139 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_140 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_141 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_142 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_143 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_144 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_145 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_146 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_147 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_148 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_149 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_150 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_151 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_152 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_153 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_154 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_155 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_156 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_157 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_158 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_159 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_160 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_161 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_162 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_163 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_164 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_165 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_166 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_167 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_168 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_169 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_170 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_171 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_172 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_173 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_174 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_175 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_176 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_177 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_178 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_179 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_180 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_181 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_182 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_183 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_184 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_185 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_186 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_187 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_188 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_189 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_190 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_191 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_192 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_193 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_194 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_195 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_196 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_197 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_198 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_199 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_200 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_201 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_202 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_203 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_204 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_205 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_206 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_207 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_208 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_209 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_210 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_211 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_212 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_213 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_214 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_215 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_216 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_217 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_218 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_219 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_220 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_221 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_222 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_223 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_224 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_225 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_226 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_227 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_228 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_229 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_230 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_231 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_232 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_233 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_234 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_235 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_236 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_237 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_238 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_239 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_240 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_241 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_242 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_243 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_244 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_245 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_246 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_247 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_248 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_249 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_250 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_251 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_252 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_253 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_254 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_255 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_256 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_257 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_258 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_259 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_260 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_261 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_262 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_263 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_264 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_265 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_266 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_267 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_268 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_269 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_270 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_271 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_272 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_273 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_274 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_275 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_276 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_277 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_278 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_279 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_280 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_281 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_282 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_283 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_284 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_285 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_286 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_287 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_288 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_289 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_290 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_291 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_292 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_293 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_294 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_295 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_296 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_297 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_298 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_299 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_300 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_301 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_302 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_303 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_304 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_305 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_306 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_307 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_308 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_309 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_310 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_311 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_312 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_313 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_314 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_315 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_316 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_317 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_318 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_319 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_320 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_321 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_322 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_323 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_324 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_325 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_326 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_327 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_328 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_329 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_330 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_331 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_332 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_333 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_334 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_335 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_336 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_337 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_338 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_339 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_340 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_341 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_342 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_343 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_344 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_345 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_346 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_347 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_348 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_349 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_350 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_351 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_352 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_353 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_354 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_355 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_356 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_357 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_358 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_359 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_360 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_361 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_362 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_363 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_364 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_365 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_366 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_367 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_368 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_369 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_370 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_371 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_372 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_373 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_374 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_375 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_376 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_377 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_378 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_379 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_380 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_381 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_382 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_383 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_384 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_385 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_386 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_387 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_388 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_389 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_390 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_391 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_392 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_393 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_394 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_395 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_396 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_397 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_398 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_399 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_400 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_401 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_402 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_403 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_404 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_405 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_406 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_407 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_408 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_409 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_410 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_411 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_412 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_413 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_414 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_415 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_416 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_417 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_418 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_419 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_420 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_421 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_422 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_423 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_424 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_425 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_426 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_427 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_428 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_429 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_430 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_431 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_432 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_433 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_434 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_435 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_436 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_437 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_438 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_439 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_440 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_441 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_442 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_443 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_444 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_445 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_446 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_447 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_448 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_449 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_450 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_451 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_452 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_453 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_454 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_455 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_456 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_457 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_458 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_459 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_460 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_461 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_462 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_463 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_464 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_465 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_466 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_467 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_468 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_469 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_470 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_471 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_472 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_473 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_474 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_475 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_476 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_477 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_478 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_479 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_480 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_481 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_482 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_483 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_484 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_485 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_486 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_487 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_488 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_489 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_490 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_491 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_492 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_493 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_494 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_495 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_496 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_497 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_498 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_499 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_500 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_501 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_502 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_503 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_504 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_505 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_506 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_507 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_508 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_509 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_510 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_511 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_512 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_513 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_514 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_515 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_516 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_517 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_518 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_519 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_520 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_521 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_522 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_523 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_524 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_525 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_526 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_527 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_528 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_529 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_530 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_531 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_532 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_533 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_534 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_535 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_536 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_537 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_538 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_539 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_540 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_541 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_542 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_543 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_544 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_545 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_546 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_547 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_548 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_549 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_550 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_551 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_552 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_553 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_554 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_555 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_556 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_557 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_558 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_559 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_560 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_561 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_562 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_563 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_564 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_565 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_566 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_567 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_568 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_569 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_570 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_571 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_572 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_573 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_574 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_575 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_576 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_577 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_578 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_579 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_580 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_581 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_582 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_583 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_584 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_585 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_586 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_587 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_588 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_589 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_590 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_591 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_592 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_593 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_594 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_595 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_596 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_597 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_598 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_599 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_600 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_601 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_602 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_603 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_604 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_605 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_606 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_607 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_608 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_609 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_610 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_611 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_612 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_613 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_614 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_615 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_616 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_617 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_618 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_619 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_620 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_621 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_622 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_623 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_624 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_625 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_626 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_627 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_628 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_629 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_630 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_631 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_632 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_633 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_634 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_635 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_636 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_637 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_638 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_639 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_640 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_641 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_642 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_643 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_644 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_645 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_646 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_647 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_648 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_649 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_650 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_651 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_652 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_653 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_654 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_655 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_656 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_657 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_658 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_659 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_660 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_661 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_662 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_663 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_664 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_665 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_666 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_667 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_668 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_669 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_670 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_671 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_672 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_673 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_674 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_675 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_676 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_677 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_678 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_679 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_680 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_681 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_682 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_683 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_684 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_685 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_686 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_687 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_688 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_689 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_690 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_691 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_692 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_693 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_694 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_695 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_696 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_697 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_698 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_699 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_700 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_701 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_702 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_703 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_704 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_705 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_706 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_707 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_708 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_709 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_710 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_711 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_712 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_713 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_714 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_715 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_716 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_717 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_718 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_719 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_720 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_721 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_722 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_723 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_724 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_725 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_726 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_727 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_728 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_729 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_730 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_731 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_732 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_733 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_734 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_735 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_736 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_737 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_738 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_739 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_740 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_741 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_742 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_743 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_744 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_745 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_746 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_747 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_748 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_749 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_750 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_751 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_752 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_753 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_754 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_755 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_756 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_757 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_758 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_759 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_760 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_761 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_762 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_763 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_764 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_765 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_766 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_767 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_768 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_769 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_770 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_771 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_772 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_773 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_774 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_775 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_776 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_777 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_778 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_779 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_780 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_781 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_782 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_783 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_784 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_785 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_786 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_787 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_788 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_789 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_790 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_791 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_792 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_793 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_794 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_795 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_796 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_797 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_798 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_799 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_800 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_801 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_802 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_803 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_804 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_805 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_806 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_807 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_808 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_809 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_810 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_811 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_812 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_813 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_814 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_815 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_816 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_817 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_818 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_819 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_820 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_821 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_822 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_823 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_824 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_825 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_826 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_827 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_828 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_829 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_830 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_831 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_832 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_833 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_834 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_835 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_836 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_837 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_838 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_839 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_840 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_841 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_842 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_843 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_844 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_845 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_846 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_847 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_848 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_849 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_850 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_851 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_852 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_853 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_854 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_855 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_856 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_857 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_858 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_859 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_860 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_861 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_862 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_863 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_864 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_865 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_866 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_867 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_868 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_869 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_870 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_871 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_872 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_873 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_874 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_875 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_876 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_877 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_878 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_879 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_880 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_881 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_882 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_883 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_884 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_885 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_886 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_887 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_888 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_889 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_890 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_891 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_892 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_893 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_894 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_895 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_896 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_897 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_898 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_899 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_900 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_901 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_902 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_903 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_904 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_905 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_906 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_907 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_908 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_909 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_910 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_911 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_912 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_913 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_914 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_915 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_916 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_917 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_918 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_919 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_920 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_921 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_922 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_923 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_924 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_925 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_926 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_927 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_928 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_929 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_930 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_931 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_932 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_933 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_934 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_935 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_936 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_937 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_938 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_939 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_940 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_941 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_942 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_943 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_944 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_945 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_946 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_947 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_948 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_949 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_950 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_951 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_952 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_953 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_954 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_955 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_956 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_957 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_958 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_959 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_960 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_961 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_962 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_963 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_964 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_965 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_966 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_967 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_968 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_969 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_970 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_971 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_972 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_973 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_974 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_975 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_976 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_977 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_978 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_979 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_980 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_981 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_982 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_983 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_984 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_985 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_986 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_987 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_988 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_989 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_990 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_991 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_992 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_993 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_994 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_995 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_996 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_997 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_998 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_999 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1000 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1001 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1002 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1003 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1004 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1005 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1006 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1007 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1008 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1009 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1010 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1011 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1012 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1013 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1014 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1015 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1016 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1017 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1018 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1019 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1020 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1021 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1022 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1023 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1024 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1025 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1026 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1027 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1028 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1029 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1030 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1031 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1032 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1033 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1034 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1035 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1036 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1037 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1038 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1039 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1040 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1041 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1042 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1043 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1044 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1045 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1046 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1047 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1048 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1049 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1050 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1051 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1052 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1053 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1054 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1055 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1056 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1057 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1058 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1059 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1060 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1061 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1062 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1063 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1064 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1065 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1066 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1067 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1068 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1069 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1070 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1071 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1072 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1073 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1074 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1075 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1076 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1077 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1078 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1079 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1080 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1081 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1082 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1083 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1084 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1085 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1086 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1087 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1088 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1089 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1090 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1091 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1092 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1093 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1094 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1095 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1096 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1097 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1098 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1099 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1100 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1101 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1102 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1103 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1104 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1105 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1106 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1107 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1108 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1109 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1110 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1111 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1112 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1113 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1114 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1115 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1116 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1117 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1118 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1119 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1120 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1121 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1122 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1123 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1124 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1125 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1126 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1127 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1128 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1129 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1130 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1131 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1132 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1133 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1134 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1135 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1136 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1137 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1138 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1139 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1140 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1141 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1142 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1143 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1144 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1145 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1146 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1147 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1148 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1149 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1150 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1151 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1152 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1153 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1154 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1155 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1156 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1157 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1158 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1159 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1160 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1161 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1162 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1163 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1164 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1165 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1166 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1167 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1168 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1169 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1170 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1171 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1172 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1173 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1174 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1175 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1176 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1177 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1178 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1179 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1180 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1181 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1182 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1183 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1184 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1185 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1186 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1187 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1188 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1189 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1190 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1191 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1192 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1193 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1194 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1195 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1196 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1197 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1198 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1199 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1200 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1201 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1202 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1203 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1204 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1205 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1206 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1207 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1208 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1209 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1210 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1211 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1212 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1213 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1214 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1215 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1216 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1217 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1218 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1219 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1220 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1221 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1222 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1223 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1224 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1225 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1226 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1227 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1228 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1229 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1230 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1231 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1232 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1233 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1234 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1235 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1236 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1237 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1238 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1239 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1240 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1241 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1242 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1243 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1244 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1245 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1246 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1247 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1248 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1249 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1250 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1251 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1252 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1253 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1254 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1255 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1256 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1257 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1258 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1259 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_1260 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_1261 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_1262 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_1263 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_1264 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_1265 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_1266 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_1267 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_1268 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_1269 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_1270 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_1271 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_1272 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_1273 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_1274 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_1275 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_1276 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_1277 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_1278 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_1279 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_1280 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_1281 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_1282 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_1283 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_1284 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_1285 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_1286 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_1287 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_1288 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_1289 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_1290 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_1291 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_1292 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_1293 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_1294 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_1295 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_1296 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_1297 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_1298 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_1299 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_1300 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_1301 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_1302 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_1303 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_1304 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_1305 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_1306 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_1307 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_1308 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_1309 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_1310 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_1311 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_1312 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_1313 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_1314 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_1315 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_1316 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_1317 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_1318 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_1319 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_1320 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_1321 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_1322 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_1323 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_1324 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_1325 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_1326 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_1327 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_1328 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_1329 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_1330 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_1331 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_1332 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_1333 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_1334 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_1335 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_1336 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_1337 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_1338 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_1339 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_1340 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_1341 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_1342 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_1343 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_1344 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_1345 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_1346 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_1347 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_1348 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_1349 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_1350 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_1351 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_1352 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_1353 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_1354 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_1355 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_1356 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_1357 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_1358 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_1359 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_1360 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_1361 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_1362 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_1363 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_1364 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_1365 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_1366 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_1367 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_1368 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_1369 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_1370 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_1371 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_1372 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_1373 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_1374 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_1375 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_1376 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_1377 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_1378 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_1379 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_1380 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_1381 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_1382 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_1383 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_1384 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_1385 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_1386 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_1387 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_1388 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_1389 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_1390 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_1391 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_1392 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_1393 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_1394 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_1395 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_1396 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_1397 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_1398 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_1399 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_1400 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_1401 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_1402 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_1403 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_1404 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_1405 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_1406 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_1407 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_1408 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_1409 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_1410 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_1411 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_1412 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_1413 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_1414 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_1415 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_1416 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_1417 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_1418 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_1419 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_1420 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_1421 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_1422 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_1423 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_1424 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_1425 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_1426 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_1427 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_1428 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_1429 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_1430 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_1431 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_1432 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_1433 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_1434 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_1435 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_1436 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_1437 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_1438 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_1439 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_1440 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_1441 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_1442 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_1443 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_1444 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_1445 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_1446 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_1447 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_1448 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_1449 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_1450 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_1451 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_1452 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_1453 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_1454 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_1455 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_1456 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_1457 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_1458 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_1459 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_1460 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_1461 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_1462 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_1463 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_1464 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_1465 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_1466 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_1467 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_1468 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_1469 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_1470 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_1471 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_1472 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_1473 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_1474 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_1475 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_1476 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_1477 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_1478 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_1479 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_1480 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_1481 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_1482 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_1483 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_1484 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_1485 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_1486 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_1487 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_1488 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_1489 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_1490 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_1491 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_1492 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_1493 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1494 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1495 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1496 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1497 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1498 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1499 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1500 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1501 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1502 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_1503 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_1504 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_1505 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_1506 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_1507 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_1508 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_1509 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_1510 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_1511 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_1512 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_1513 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_1514 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_1515 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_1516 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_1517 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_1518 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_1519 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_1520 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_1521 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_1522 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_1523 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_1524 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_1525 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_1526 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_1527 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_1528 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_1529 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_1530 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_1531 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_1532 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_1533 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_1534 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_1535 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_1536 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_1537 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_1538 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_1539 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_1540 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_1541 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_1542 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_1543 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_1544 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_1545 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_1546 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_1547 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_1548 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_1549 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_1550 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_1551 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_1552 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_1553 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_1554 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_1555 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_1556 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_1557 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_1558 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_1559 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_1560 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_1561 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_1562 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_1563 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_1564 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_1565 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_1566 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_1567 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_1568 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_1569 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_1570 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_1571 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_1572 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_1573 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_1574 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1575 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1576 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1577 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1578 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1579 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1580 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1581 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1582 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1583 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_1584 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_1585 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_1586 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_1587 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_1588 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_1589 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_1590 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_1591 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_1592 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_1593 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_1594 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_1595 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_1596 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_1597 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_1598 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_1599 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_1600 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_1601 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_1602 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_1603 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_1604 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_1605 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_1606 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_1607 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_1608 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_1609 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_1610 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_1611 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_1612 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_1613 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_1614 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_1615 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_1616 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_1617 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_1618 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_1619 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_1620 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_1621 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_1622 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_1623 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_1624 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_1625 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_1626 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_1627 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_1628 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_1629 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_1630 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_1631 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_1632 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_1633 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_1634 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_1635 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_1636 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_1637 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_1638 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_1639 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_1640 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_1641 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_1642 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_1643 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_1644 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_1645 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_1646 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_1647 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_1648 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_1649 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_1650 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_1651 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_1652 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_1653 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_1654 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_1655 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_1656 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_1657 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_1658 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_1659 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_1660 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_1661 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_1662 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_1663 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_1664 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_1665 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_1666 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_1667 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_1668 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_1669 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_1670 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_1671 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_1672 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_1673 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_1674 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_1675 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_1676 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_1677 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_1678 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_1679 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_1680 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_1681 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_1682 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_1683 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_1684 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_1685 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_1686 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_1687 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_1688 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_1689 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_1690 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_1691 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_1692 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_1693 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_1694 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_1695 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_1696 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_1697 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_1698 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_1699 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_1700 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_1701 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_1702 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_1703 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_1704 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_1705 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_1706 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_1707 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_1708 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_1709 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_1710 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_1711 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_1712 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_1713 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_1714 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_1715 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_1716 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_1717 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_1718 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_1719 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_1720 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_1721 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_1722 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_1723 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_1724 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_1725 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_1726 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_1727 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_1728 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_1729 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_1730 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_1731 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_1732 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_1733 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_1734 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_1735 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_1736 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_1737 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_1738 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_1739 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_1740 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_1741 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_1742 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_1743 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_1744 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_1745 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_1746 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_1747 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_1748 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_1749 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_1750 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_1751 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_1752 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_1753 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_1754 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_1755 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_1756 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_1757 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_1758 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_1759 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_1760 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_1761 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_1762 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_1763 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_1764 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_1765 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_1766 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_1767 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_1768 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_1769 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_1770 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_1771 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_1772 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_1773 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_1774 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_1775 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_1776 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_1777 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_1778 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_1779 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_1780 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_1781 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_1782 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_1783 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_1784 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_1785 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_1786 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_1787 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_1788 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_1789 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_1790 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_1791 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_1792 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_1793 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_1794 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_1795 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_1796 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_1797 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_1798 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_1799 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_1800 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_1801 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_1802 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_1803 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_1804 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_1805 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_1806 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_1807 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_1808 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_1809 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_1810 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_1811 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_1812 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_1813 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_1814 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_1815 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_1816 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_1817 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_1818 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_1819 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_1820 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_1821 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_1822 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_1823 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_1824 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_1825 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_1826 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_1827 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_1828 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_1829 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_1830 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_1831 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_1832 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_1833 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_1834 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_1835 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_1836 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_1837 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_1838 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_1839 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_1840 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_1841 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_1842 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_1843 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_1844 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_1845 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_1846 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_1847 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_1848 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_1849 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_1850 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_1851 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_1852 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_1853 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_1854 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_1855 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_1856 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_1857 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_1858 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_1859 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_1860 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_1861 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_1862 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_1863 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_1864 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_1865 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_1866 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_1867 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_1868 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_1869 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_1870 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_1871 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_1872 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_1873 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_1874 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_1875 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_1876 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_1877 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_1878 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_1879 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_1880 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_1881 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_1882 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_1883 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_1884 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_1885 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_1886 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_1887 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_1888 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_1889 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_1890 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_1891 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_1892 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_1893 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_1894 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_1895 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_1896 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_1897 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_1898 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_1899 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_1900 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_1901 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_1902 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_1903 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_1904 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_1905 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_1906 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_1907 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_1908 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_1909 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_1910 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_1911 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_1912 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_1913 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_1914 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_1915 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_1916 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_1917 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_1918 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_1919 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_1920 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_1921 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_1922 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_1923 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_1924 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_1925 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_1926 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_1927 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_1928 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_1929 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_1930 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_1931 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_1932 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_1933 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_1934 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_1935 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_1936 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_1937 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_1938 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_1939 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_1940 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_1941 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_1942 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_1943 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_1944 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_1945 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_1946 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_1947 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_1948 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_1949 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_1950 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_1951 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_1952 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_1953 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_1954 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_1955 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_1956 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_1957 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_1958 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_1959 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_1960 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_1961 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_1962 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_1963 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_1964 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_1965 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_1966 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_1967 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_1968 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_1969 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_1970 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_1971 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_1972 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_1973 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_1974 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_1975 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_1976 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_1977 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_1978 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_1979 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_1980 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_1981 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_1982 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_1983 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_1984 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_1985 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_1986 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_1987 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_1988 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_1989 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_1990 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_1991 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_1992 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_1993 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_1994 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_1995 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_1996 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_1997 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_1998 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_1999 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_2000 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_2001 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_2002 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_2003 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_2004 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_2005 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_2006 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_2007 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_2008 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_2009 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_2010 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_2011 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_2012 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_2013 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_2014 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_2015 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_2016 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_2017 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_2018 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_2019 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_2020 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_2021 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_2022 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_2023 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_2024 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_2025 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_2026 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_2027 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_2028 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_2029 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_2030 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_2031 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_2032 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_2033 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_2034 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_2035 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_2036 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_2037 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_2038 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_2039 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_2040 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_2041 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_2042 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_2043 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_2044 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_2045 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_2046 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_2047 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_2048 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_2049 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_2050 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_2051 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_2052 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_2053 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_2054 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_2055 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_2056 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_2057 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_2058 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_2059 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_2060 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_2061 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_2062 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_2063 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_2064 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_2065 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_2066 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_2067 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_2068 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_2069 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_2070 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_2071 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_2072 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_2073 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_2074 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_2075 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_2076 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_2077 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_2078 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_2079 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_2080 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_2081 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_2082 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_2083 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_2084 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_2085 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_2086 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_2087 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_2088 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_2089 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_2090 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_2091 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_2092 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_2093 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_2094 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_2095 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_2096 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_2097 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_2098 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_2099 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_2100 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_2101 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_2102 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_2103 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_2104 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_2105 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_2106 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_2107 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_2108 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_2109 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_2110 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_2111 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_2112 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_2113 ();
 sky130_fd_sc_hs__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_2114 ();
 sky130_fd_sc_hs__buf_4 wire9 (.A(net11),
    .X(net9));
 sky130_fd_sc_hs__buf_4 load_slew10 (.A(net11),
    .X(net212));
 sky130_fd_sc_hs__buf_4 load_slew11 (.A(net10),
    .X(net11));
 sky130_fd_sc_hs__buf_8 wire12 (.A(net211),
    .X(net12));
 sky130_fd_sc_hs__buf_8 load_slew13 (.A(net14),
    .X(net13));
 sky130_fd_sc_hs__buf_8 max_cap14 (.A(net14),
    .X(net207));
 sky130_fd_sc_hs__buf_8 load_slew15 (.A(net15),
    .X(net197));
 sky130_fd_sc_hs__buf_8 wire16 (.A(net16),
    .X(net196));
 sky130_fd_sc_hs__dlygate4sd1_1 input1 (.A(alu_instr_first_cycle_i),
    .X(net1));
 sky130_fd_sc_hs__dlygate4sd1_1 input2 (.A(alu_operand_a_i[0]),
    .X(net2));
 sky130_fd_sc_hs__dlygate4sd1_1 input3 (.A(alu_operand_a_i[10]),
    .X(net3));
 sky130_fd_sc_hs__dlygate4sd1_1 input4 (.A(alu_operand_a_i[11]),
    .X(net4));
 sky130_fd_sc_hs__dlygate4sd1_1 input5 (.A(alu_operand_a_i[12]),
    .X(net5));
 sky130_fd_sc_hs__dlygate4sd1_1 input6 (.A(alu_operand_a_i[13]),
    .X(net6));
 sky130_fd_sc_hs__dlygate4sd1_1 input7 (.A(alu_operand_a_i[14]),
    .X(net7));
 sky130_fd_sc_hs__dlygate4sd1_1 input8 (.A(alu_operand_a_i[15]),
    .X(net8));
 sky130_fd_sc_hs__dlygate4sd1_1 input9 (.A(alu_operand_a_i[16]),
    .X(net17));
 sky130_fd_sc_hs__dlygate4sd1_1 input10 (.A(alu_operand_a_i[17]),
    .X(net18));
 sky130_fd_sc_hs__dlygate4sd1_1 input11 (.A(alu_operand_a_i[18]),
    .X(net19));
 sky130_fd_sc_hs__dlygate4sd1_1 input12 (.A(alu_operand_a_i[19]),
    .X(net20));
 sky130_fd_sc_hs__dlygate4sd1_1 input13 (.A(alu_operand_a_i[1]),
    .X(net21));
 sky130_fd_sc_hs__dlygate4sd1_1 input14 (.A(alu_operand_a_i[20]),
    .X(net22));
 sky130_fd_sc_hs__dlygate4sd1_1 input15 (.A(alu_operand_a_i[21]),
    .X(net23));
 sky130_fd_sc_hs__dlygate4sd1_1 input16 (.A(alu_operand_a_i[22]),
    .X(net24));
 sky130_fd_sc_hs__dlygate4sd1_1 input17 (.A(alu_operand_a_i[23]),
    .X(net25));
 sky130_fd_sc_hs__dlygate4sd1_1 input18 (.A(alu_operand_a_i[24]),
    .X(net26));
 sky130_fd_sc_hs__dlygate4sd1_1 input19 (.A(alu_operand_a_i[25]),
    .X(net27));
 sky130_fd_sc_hs__dlygate4sd1_1 input20 (.A(alu_operand_a_i[26]),
    .X(net28));
 sky130_fd_sc_hs__dlygate4sd1_1 input21 (.A(alu_operand_a_i[27]),
    .X(net29));
 sky130_fd_sc_hs__dlygate4sd1_1 input22 (.A(alu_operand_a_i[28]),
    .X(net30));
 sky130_fd_sc_hs__dlygate4sd1_1 input23 (.A(alu_operand_a_i[29]),
    .X(net31));
 sky130_fd_sc_hs__dlygate4sd1_1 input24 (.A(alu_operand_a_i[2]),
    .X(net32));
 sky130_fd_sc_hs__dlygate4sd1_1 input25 (.A(alu_operand_a_i[30]),
    .X(net33));
 sky130_fd_sc_hs__dlygate4sd1_1 input26 (.A(alu_operand_a_i[31]),
    .X(net34));
 sky130_fd_sc_hs__dlygate4sd1_1 input27 (.A(alu_operand_a_i[3]),
    .X(net35));
 sky130_fd_sc_hs__dlygate4sd1_1 input28 (.A(alu_operand_a_i[4]),
    .X(net36));
 sky130_fd_sc_hs__dlygate4sd1_1 input29 (.A(alu_operand_a_i[5]),
    .X(net37));
 sky130_fd_sc_hs__dlygate4sd1_1 input30 (.A(alu_operand_a_i[6]),
    .X(net38));
 sky130_fd_sc_hs__dlygate4sd1_1 input31 (.A(alu_operand_a_i[7]),
    .X(net39));
 sky130_fd_sc_hs__dlygate4sd1_1 input32 (.A(alu_operand_a_i[8]),
    .X(net40));
 sky130_fd_sc_hs__dlygate4sd1_1 input33 (.A(alu_operand_a_i[9]),
    .X(net41));
 sky130_fd_sc_hs__dlygate4sd1_1 input34 (.A(alu_operand_b_i[0]),
    .X(net42));
 sky130_fd_sc_hs__dlygate4sd1_1 input35 (.A(alu_operand_b_i[10]),
    .X(net43));
 sky130_fd_sc_hs__dlygate4sd1_1 input36 (.A(alu_operand_b_i[11]),
    .X(net44));
 sky130_fd_sc_hs__dlygate4sd1_1 input37 (.A(alu_operand_b_i[12]),
    .X(net45));
 sky130_fd_sc_hs__dlygate4sd1_1 input38 (.A(alu_operand_b_i[13]),
    .X(net46));
 sky130_fd_sc_hs__dlygate4sd1_1 input39 (.A(alu_operand_b_i[14]),
    .X(net47));
 sky130_fd_sc_hs__dlygate4sd1_1 input40 (.A(alu_operand_b_i[15]),
    .X(net48));
 sky130_fd_sc_hs__dlygate4sd1_1 input41 (.A(alu_operand_b_i[16]),
    .X(net49));
 sky130_fd_sc_hs__dlygate4sd1_1 input42 (.A(alu_operand_b_i[17]),
    .X(net50));
 sky130_fd_sc_hs__dlygate4sd1_1 input43 (.A(alu_operand_b_i[18]),
    .X(net51));
 sky130_fd_sc_hs__dlygate4sd1_1 input44 (.A(alu_operand_b_i[19]),
    .X(net52));
 sky130_fd_sc_hs__dlygate4sd1_1 input45 (.A(alu_operand_b_i[1]),
    .X(net53));
 sky130_fd_sc_hs__dlygate4sd1_1 input46 (.A(alu_operand_b_i[20]),
    .X(net54));
 sky130_fd_sc_hs__dlygate4sd1_1 input47 (.A(alu_operand_b_i[21]),
    .X(net55));
 sky130_fd_sc_hs__dlygate4sd1_1 input48 (.A(alu_operand_b_i[22]),
    .X(net56));
 sky130_fd_sc_hs__dlygate4sd1_1 input49 (.A(alu_operand_b_i[23]),
    .X(net57));
 sky130_fd_sc_hs__dlygate4sd1_1 input50 (.A(alu_operand_b_i[24]),
    .X(net58));
 sky130_fd_sc_hs__dlygate4sd1_1 input51 (.A(alu_operand_b_i[25]),
    .X(net59));
 sky130_fd_sc_hs__dlygate4sd1_1 input52 (.A(alu_operand_b_i[26]),
    .X(net60));
 sky130_fd_sc_hs__dlygate4sd1_1 input53 (.A(alu_operand_b_i[27]),
    .X(net61));
 sky130_fd_sc_hs__dlygate4sd1_1 input54 (.A(alu_operand_b_i[28]),
    .X(net62));
 sky130_fd_sc_hs__dlygate4sd1_1 input55 (.A(alu_operand_b_i[29]),
    .X(net63));
 sky130_fd_sc_hs__dlygate4sd1_1 input56 (.A(alu_operand_b_i[2]),
    .X(net64));
 sky130_fd_sc_hs__dlygate4sd1_1 input57 (.A(alu_operand_b_i[30]),
    .X(net65));
 sky130_fd_sc_hs__dlygate4sd1_1 input58 (.A(alu_operand_b_i[31]),
    .X(net66));
 sky130_fd_sc_hs__dlygate4sd1_1 input59 (.A(alu_operand_b_i[3]),
    .X(net67));
 sky130_fd_sc_hs__dlygate4sd1_1 input60 (.A(alu_operand_b_i[4]),
    .X(net68));
 sky130_fd_sc_hs__dlygate4sd1_1 input61 (.A(alu_operand_b_i[5]),
    .X(net69));
 sky130_fd_sc_hs__dlygate4sd1_1 input62 (.A(alu_operand_b_i[6]),
    .X(net70));
 sky130_fd_sc_hs__dlygate4sd1_1 input63 (.A(alu_operand_b_i[7]),
    .X(net71));
 sky130_fd_sc_hs__dlygate4sd1_1 input64 (.A(alu_operand_b_i[8]),
    .X(net72));
 sky130_fd_sc_hs__dlygate4sd1_1 input65 (.A(alu_operand_b_i[9]),
    .X(net73));
 sky130_fd_sc_hs__dlygate4sd1_1 input66 (.A(alu_operator_i[0]),
    .X(net74));
 sky130_fd_sc_hs__dlygate4sd1_1 input67 (.A(alu_operator_i[1]),
    .X(net75));
 sky130_fd_sc_hs__dlygate4sd1_1 input68 (.A(alu_operator_i[4]),
    .X(net76));
 sky130_fd_sc_hs__dlygate4sd1_1 input69 (.A(alu_operator_i[5]),
    .X(net77));
 sky130_fd_sc_hs__dlygate4sd1_1 input70 (.A(data_ind_timing_i),
    .X(net78));
 sky130_fd_sc_hs__dlygate4sd1_1 input71 (.A(div_en_i),
    .X(net79));
 sky130_fd_sc_hs__dlygate4sd1_1 input72 (.A(div_sel_i),
    .X(net80));
 sky130_fd_sc_hs__dlygate4sd1_1 input73 (.A(imd_val_q_i[0]),
    .X(net81));
 sky130_fd_sc_hs__dlygate4sd1_1 input74 (.A(imd_val_q_i[10]),
    .X(net82));
 sky130_fd_sc_hs__dlygate4sd1_1 input75 (.A(imd_val_q_i[11]),
    .X(net83));
 sky130_fd_sc_hs__dlygate4sd1_1 input76 (.A(imd_val_q_i[12]),
    .X(net84));
 sky130_fd_sc_hs__dlygate4sd1_1 input77 (.A(imd_val_q_i[13]),
    .X(net85));
 sky130_fd_sc_hs__dlygate4sd1_1 input78 (.A(imd_val_q_i[14]),
    .X(net86));
 sky130_fd_sc_hs__dlygate4sd1_1 input79 (.A(imd_val_q_i[15]),
    .X(net87));
 sky130_fd_sc_hs__dlygate4sd1_1 input80 (.A(imd_val_q_i[16]),
    .X(net88));
 sky130_fd_sc_hs__dlygate4sd1_1 input81 (.A(imd_val_q_i[17]),
    .X(net89));
 sky130_fd_sc_hs__dlygate4sd1_1 input82 (.A(imd_val_q_i[18]),
    .X(net90));
 sky130_fd_sc_hs__dlygate4sd1_1 input83 (.A(imd_val_q_i[19]),
    .X(net91));
 sky130_fd_sc_hs__dlygate4sd1_1 input84 (.A(imd_val_q_i[1]),
    .X(net92));
 sky130_fd_sc_hs__dlygate4sd1_1 input85 (.A(imd_val_q_i[20]),
    .X(net93));
 sky130_fd_sc_hs__dlygate4sd1_1 input86 (.A(imd_val_q_i[21]),
    .X(net94));
 sky130_fd_sc_hs__dlygate4sd1_1 input87 (.A(imd_val_q_i[22]),
    .X(net95));
 sky130_fd_sc_hs__dlygate4sd1_1 input88 (.A(imd_val_q_i[23]),
    .X(net96));
 sky130_fd_sc_hs__dlygate4sd1_1 input89 (.A(imd_val_q_i[24]),
    .X(net97));
 sky130_fd_sc_hs__dlygate4sd1_1 input90 (.A(imd_val_q_i[25]),
    .X(net98));
 sky130_fd_sc_hs__dlygate4sd1_1 input91 (.A(imd_val_q_i[26]),
    .X(net99));
 sky130_fd_sc_hs__dlygate4sd1_1 input92 (.A(imd_val_q_i[27]),
    .X(net100));
 sky130_fd_sc_hs__dlygate4sd1_1 input93 (.A(imd_val_q_i[28]),
    .X(net101));
 sky130_fd_sc_hs__dlygate4sd1_1 input94 (.A(imd_val_q_i[29]),
    .X(net102));
 sky130_fd_sc_hs__dlygate4sd1_1 input95 (.A(imd_val_q_i[2]),
    .X(net103));
 sky130_fd_sc_hs__dlygate4sd1_1 input96 (.A(imd_val_q_i[30]),
    .X(net104));
 sky130_fd_sc_hs__dlygate4sd1_1 input97 (.A(imd_val_q_i[31]),
    .X(net105));
 sky130_fd_sc_hs__dlygate4sd1_1 input98 (.A(imd_val_q_i[3]),
    .X(net106));
 sky130_fd_sc_hs__dlygate4sd1_1 input99 (.A(imd_val_q_i[49]),
    .X(net107));
 sky130_fd_sc_hs__dlygate4sd1_1 input100 (.A(imd_val_q_i[4]),
    .X(net108));
 sky130_fd_sc_hs__buf_16 input101 (.A(imd_val_q_i[55]),
    .X(net109));
 sky130_fd_sc_hs__dlygate4sd1_1 input102 (.A(imd_val_q_i[5]),
    .X(net110));
 sky130_fd_sc_hs__dlygate4sd1_1 input103 (.A(imd_val_q_i[62]),
    .X(net111));
 sky130_fd_sc_hs__dlygate4sd1_1 input104 (.A(imd_val_q_i[63]),
    .X(net112));
 sky130_fd_sc_hs__dlygate4sd1_1 input105 (.A(imd_val_q_i[65]),
    .X(net113));
 sky130_fd_sc_hs__dlygate4sd1_1 input106 (.A(imd_val_q_i[66]),
    .X(net114));
 sky130_fd_sc_hs__dlygate4sd1_1 input107 (.A(imd_val_q_i[67]),
    .X(net115));
 sky130_fd_sc_hs__dlygate4sd1_1 input108 (.A(imd_val_q_i[6]),
    .X(net116));
 sky130_fd_sc_hs__dlygate4sd1_1 input109 (.A(imd_val_q_i[7]),
    .X(net117));
 sky130_fd_sc_hs__dlygate4sd1_1 input110 (.A(imd_val_q_i[8]),
    .X(net118));
 sky130_fd_sc_hs__dlygate4sd1_1 input111 (.A(imd_val_q_i[9]),
    .X(net119));
 sky130_fd_sc_hs__dlygate4sd1_1 input112 (.A(mult_en_i),
    .X(net120));
 sky130_fd_sc_hs__dlygate4sd1_1 input113 (.A(multdiv_operand_a_i[0]),
    .X(net121));
 sky130_fd_sc_hs__dlygate4sd1_1 input114 (.A(multdiv_operand_a_i[10]),
    .X(net122));
 sky130_fd_sc_hs__dlygate4sd1_1 input115 (.A(multdiv_operand_a_i[11]),
    .X(net123));
 sky130_fd_sc_hs__dlygate4sd1_1 input116 (.A(multdiv_operand_a_i[12]),
    .X(net124));
 sky130_fd_sc_hs__dlygate4sd1_1 input117 (.A(multdiv_operand_a_i[13]),
    .X(net125));
 sky130_fd_sc_hs__dlygate4sd1_1 input118 (.A(multdiv_operand_a_i[14]),
    .X(net126));
 sky130_fd_sc_hs__dlygate4sd1_1 input119 (.A(multdiv_operand_a_i[15]),
    .X(net127));
 sky130_fd_sc_hs__dlygate4sd1_1 input120 (.A(multdiv_operand_a_i[16]),
    .X(net128));
 sky130_fd_sc_hs__dlygate4sd1_1 input121 (.A(multdiv_operand_a_i[17]),
    .X(net129));
 sky130_fd_sc_hs__dlygate4sd1_1 input122 (.A(multdiv_operand_a_i[18]),
    .X(net130));
 sky130_fd_sc_hs__dlygate4sd1_1 input123 (.A(multdiv_operand_a_i[19]),
    .X(net131));
 sky130_fd_sc_hs__dlygate4sd1_1 input124 (.A(multdiv_operand_a_i[1]),
    .X(net132));
 sky130_fd_sc_hs__dlygate4sd1_1 input125 (.A(multdiv_operand_a_i[20]),
    .X(net133));
 sky130_fd_sc_hs__dlygate4sd1_1 input126 (.A(multdiv_operand_a_i[21]),
    .X(net134));
 sky130_fd_sc_hs__dlygate4sd1_1 input127 (.A(multdiv_operand_a_i[22]),
    .X(net135));
 sky130_fd_sc_hs__dlygate4sd1_1 input128 (.A(multdiv_operand_a_i[23]),
    .X(net136));
 sky130_fd_sc_hs__dlygate4sd1_1 input129 (.A(multdiv_operand_a_i[24]),
    .X(net137));
 sky130_fd_sc_hs__dlygate4sd1_1 input130 (.A(multdiv_operand_a_i[25]),
    .X(net138));
 sky130_fd_sc_hs__dlygate4sd1_1 input131 (.A(multdiv_operand_a_i[26]),
    .X(net139));
 sky130_fd_sc_hs__dlygate4sd1_1 input132 (.A(multdiv_operand_a_i[27]),
    .X(net140));
 sky130_fd_sc_hs__dlygate4sd1_1 input133 (.A(multdiv_operand_a_i[28]),
    .X(net141));
 sky130_fd_sc_hs__dlygate4sd1_1 input134 (.A(multdiv_operand_a_i[29]),
    .X(net142));
 sky130_fd_sc_hs__dlygate4sd1_1 input135 (.A(multdiv_operand_a_i[2]),
    .X(net143));
 sky130_fd_sc_hs__dlygate4sd1_1 input136 (.A(multdiv_operand_a_i[30]),
    .X(net144));
 sky130_fd_sc_hs__dlygate4sd1_1 input137 (.A(multdiv_operand_a_i[31]),
    .X(net145));
 sky130_fd_sc_hs__dlygate4sd1_1 input138 (.A(multdiv_operand_a_i[3]),
    .X(net146));
 sky130_fd_sc_hs__dlygate4sd1_1 input139 (.A(multdiv_operand_a_i[4]),
    .X(net147));
 sky130_fd_sc_hs__dlygate4sd1_1 input140 (.A(multdiv_operand_a_i[5]),
    .X(net148));
 sky130_fd_sc_hs__dlygate4sd1_1 input141 (.A(multdiv_operand_a_i[6]),
    .X(net149));
 sky130_fd_sc_hs__dlygate4sd1_1 input142 (.A(multdiv_operand_a_i[7]),
    .X(net150));
 sky130_fd_sc_hs__dlygate4sd1_1 input143 (.A(multdiv_operand_a_i[8]),
    .X(net151));
 sky130_fd_sc_hs__dlygate4sd1_1 input144 (.A(multdiv_operand_a_i[9]),
    .X(net152));
 sky130_fd_sc_hs__dlygate4sd1_1 input145 (.A(multdiv_operand_b_i[0]),
    .X(net153));
 sky130_fd_sc_hs__dlygate4sd1_1 input146 (.A(multdiv_operand_b_i[10]),
    .X(net154));
 sky130_fd_sc_hs__dlygate4sd1_1 input147 (.A(multdiv_operand_b_i[11]),
    .X(net155));
 sky130_fd_sc_hs__dlygate4sd1_1 input148 (.A(multdiv_operand_b_i[12]),
    .X(net156));
 sky130_fd_sc_hs__dlygate4sd1_1 input149 (.A(multdiv_operand_b_i[13]),
    .X(net157));
 sky130_fd_sc_hs__dlygate4sd1_1 input150 (.A(multdiv_operand_b_i[14]),
    .X(net158));
 sky130_fd_sc_hs__dlygate4sd1_1 input151 (.A(multdiv_operand_b_i[15]),
    .X(net159));
 sky130_fd_sc_hs__dlygate4sd1_1 input152 (.A(multdiv_operand_b_i[16]),
    .X(net160));
 sky130_fd_sc_hs__dlygate4sd1_1 input153 (.A(multdiv_operand_b_i[17]),
    .X(net161));
 sky130_fd_sc_hs__dlygate4sd1_1 input154 (.A(multdiv_operand_b_i[18]),
    .X(net162));
 sky130_fd_sc_hs__dlygate4sd1_1 input155 (.A(multdiv_operand_b_i[19]),
    .X(net163));
 sky130_fd_sc_hs__dlygate4sd1_1 input156 (.A(multdiv_operand_b_i[1]),
    .X(net164));
 sky130_fd_sc_hs__dlygate4sd1_1 input157 (.A(multdiv_operand_b_i[20]),
    .X(net165));
 sky130_fd_sc_hs__dlygate4sd1_1 input158 (.A(multdiv_operand_b_i[21]),
    .X(net166));
 sky130_fd_sc_hs__dlygate4sd1_1 input159 (.A(multdiv_operand_b_i[22]),
    .X(net167));
 sky130_fd_sc_hs__dlygate4sd1_1 input160 (.A(multdiv_operand_b_i[23]),
    .X(net168));
 sky130_fd_sc_hs__dlygate4sd1_1 input161 (.A(multdiv_operand_b_i[24]),
    .X(net169));
 sky130_fd_sc_hs__dlygate4sd1_1 input162 (.A(multdiv_operand_b_i[25]),
    .X(net170));
 sky130_fd_sc_hs__dlygate4sd1_1 input163 (.A(multdiv_operand_b_i[26]),
    .X(net171));
 sky130_fd_sc_hs__dlygate4sd1_1 input164 (.A(multdiv_operand_b_i[27]),
    .X(net172));
 sky130_fd_sc_hs__dlygate4sd1_1 input165 (.A(multdiv_operand_b_i[28]),
    .X(net173));
 sky130_fd_sc_hs__dlygate4sd1_1 input166 (.A(multdiv_operand_b_i[29]),
    .X(net174));
 sky130_fd_sc_hs__dlygate4sd1_1 input167 (.A(multdiv_operand_b_i[2]),
    .X(net175));
 sky130_fd_sc_hs__dlygate4sd1_1 input168 (.A(multdiv_operand_b_i[30]),
    .X(net176));
 sky130_fd_sc_hs__dlygate4sd1_1 input169 (.A(multdiv_operand_b_i[31]),
    .X(net177));
 sky130_fd_sc_hs__dlygate4sd1_1 input170 (.A(multdiv_operand_b_i[3]),
    .X(net178));
 sky130_fd_sc_hs__dlygate4sd1_1 input171 (.A(multdiv_operand_b_i[4]),
    .X(net179));
 sky130_fd_sc_hs__dlygate4sd1_1 input172 (.A(multdiv_operand_b_i[5]),
    .X(net180));
 sky130_fd_sc_hs__dlygate4sd1_1 input173 (.A(multdiv_operand_b_i[6]),
    .X(net181));
 sky130_fd_sc_hs__dlygate4sd1_1 input174 (.A(multdiv_operand_b_i[7]),
    .X(net182));
 sky130_fd_sc_hs__dlygate4sd1_1 input175 (.A(multdiv_operand_b_i[8]),
    .X(net183));
 sky130_fd_sc_hs__dlygate4sd1_1 input176 (.A(multdiv_operand_b_i[9]),
    .X(net184));
 sky130_fd_sc_hs__dlygate4sd1_1 input177 (.A(multdiv_operator_i[0]),
    .X(net185));
 sky130_fd_sc_hs__dlygate4sd1_1 input178 (.A(multdiv_operator_i[1]),
    .X(net186));
 sky130_fd_sc_hs__dlygate4sd1_1 input179 (.A(multdiv_ready_id_i),
    .X(net187));
 sky130_fd_sc_hs__dlygate4sd1_1 input180 (.A(multdiv_signed_mode_i[0]),
    .X(net188));
 sky130_fd_sc_hs__dlygate4sd1_1 input181 (.A(multdiv_signed_mode_i[1]),
    .X(net189));
 sky130_fd_sc_hs__dlygate4sd1_1 input182 (.A(rst_ni),
    .X(net190));
 sky130_fd_sc_hs__dlygate4sd1_1 output183 (.A(net191),
    .X(alu_adder_result_ex_o[0]));
 sky130_fd_sc_hs__dlygate4sd1_1 output184 (.A(net192),
    .X(alu_adder_result_ex_o[10]));
 sky130_fd_sc_hs__dlygate4sd1_1 output185 (.A(net365),
    .X(alu_adder_result_ex_o[11]));
 sky130_fd_sc_hs__dlygate4sd1_1 output186 (.A(net194),
    .X(alu_adder_result_ex_o[12]));
 sky130_fd_sc_hs__dlygate4sd1_1 output187 (.A(net195),
    .X(alu_adder_result_ex_o[13]));
 sky130_fd_sc_hs__dlygate4sd1_1 output188 (.A(net196),
    .X(alu_adder_result_ex_o[14]));
 sky130_fd_sc_hs__dlygate4sd1_1 output189 (.A(net197),
    .X(alu_adder_result_ex_o[15]));
 sky130_fd_sc_hs__dlygate4sd1_1 output190 (.A(net198),
    .X(alu_adder_result_ex_o[16]));
 sky130_fd_sc_hs__dlygate4sd1_1 output191 (.A(net199),
    .X(alu_adder_result_ex_o[17]));
 sky130_fd_sc_hs__dlygate4sd1_1 output192 (.A(net200),
    .X(alu_adder_result_ex_o[18]));
 sky130_fd_sc_hs__dlygate4sd1_1 output193 (.A(net201),
    .X(alu_adder_result_ex_o[19]));
 sky130_fd_sc_hs__dlygate4sd1_1 output194 (.A(net202),
    .X(alu_adder_result_ex_o[1]));
 sky130_fd_sc_hs__dlygate4sd1_1 output195 (.A(net203),
    .X(alu_adder_result_ex_o[20]));
 sky130_fd_sc_hs__dlygate4sd1_1 output196 (.A(net204),
    .X(alu_adder_result_ex_o[21]));
 sky130_fd_sc_hs__dlygate4sd1_1 output197 (.A(net205),
    .X(alu_adder_result_ex_o[22]));
 sky130_fd_sc_hs__dlygate4sd1_1 output198 (.A(net206),
    .X(alu_adder_result_ex_o[23]));
 sky130_fd_sc_hs__dlygate4sd1_1 output199 (.A(net207),
    .X(alu_adder_result_ex_o[24]));
 sky130_fd_sc_hs__dlygate4sd1_1 output200 (.A(net208),
    .X(alu_adder_result_ex_o[25]));
 sky130_fd_sc_hs__dlygate4sd1_1 output201 (.A(net209),
    .X(alu_adder_result_ex_o[26]));
 sky130_fd_sc_hs__dlygate4sd1_1 output202 (.A(net210),
    .X(alu_adder_result_ex_o[27]));
 sky130_fd_sc_hs__dlygate4sd1_1 output203 (.A(net211),
    .X(alu_adder_result_ex_o[28]));
 sky130_fd_sc_hs__dlygate4sd1_1 output204 (.A(net212),
    .X(alu_adder_result_ex_o[29]));
 sky130_fd_sc_hs__dlygate4sd1_1 output205 (.A(net213),
    .X(alu_adder_result_ex_o[2]));
 sky130_fd_sc_hs__dlygate4sd1_1 output206 (.A(net214),
    .X(alu_adder_result_ex_o[30]));
 sky130_fd_sc_hs__dlygate4sd1_1 output207 (.A(net215),
    .X(alu_adder_result_ex_o[31]));
 sky130_fd_sc_hs__dlygate4sd1_1 output208 (.A(net216),
    .X(alu_adder_result_ex_o[3]));
 sky130_fd_sc_hs__dlygate4sd1_1 output209 (.A(net217),
    .X(alu_adder_result_ex_o[4]));
 sky130_fd_sc_hs__dlygate4sd1_1 output210 (.A(net218),
    .X(alu_adder_result_ex_o[5]));
 sky130_fd_sc_hs__dlygate4sd1_1 output211 (.A(net219),
    .X(alu_adder_result_ex_o[6]));
 sky130_fd_sc_hs__dlygate4sd1_1 output212 (.A(net220),
    .X(alu_adder_result_ex_o[7]));
 sky130_fd_sc_hs__dlygate4sd1_1 output213 (.A(net221),
    .X(alu_adder_result_ex_o[8]));
 sky130_fd_sc_hs__dlygate4sd1_1 output214 (.A(net222),
    .X(alu_adder_result_ex_o[9]));
 sky130_fd_sc_hs__dlygate4sd1_1 output215 (.A(net223),
    .X(branch_decision_o));
 sky130_fd_sc_hs__dlygate4sd1_1 output216 (.A(net224),
    .X(branch_target_o[0]));
 sky130_fd_sc_hs__dlygate4sd1_1 output217 (.A(net225),
    .X(branch_target_o[10]));
 sky130_fd_sc_hs__dlygate4sd1_1 output218 (.A(net226),
    .X(branch_target_o[11]));
 sky130_fd_sc_hs__dlygate4sd1_1 output219 (.A(net227),
    .X(branch_target_o[12]));
 sky130_fd_sc_hs__dlygate4sd1_1 output220 (.A(net228),
    .X(branch_target_o[13]));
 sky130_fd_sc_hs__dlygate4sd1_1 output221 (.A(net229),
    .X(branch_target_o[14]));
 sky130_fd_sc_hs__dlygate4sd1_1 output222 (.A(net230),
    .X(branch_target_o[15]));
 sky130_fd_sc_hs__dlygate4sd1_1 output223 (.A(net231),
    .X(branch_target_o[16]));
 sky130_fd_sc_hs__dlygate4sd1_1 output224 (.A(net232),
    .X(branch_target_o[17]));
 sky130_fd_sc_hs__dlygate4sd1_1 output225 (.A(net233),
    .X(branch_target_o[18]));
 sky130_fd_sc_hs__dlygate4sd1_1 output226 (.A(net234),
    .X(branch_target_o[19]));
 sky130_fd_sc_hs__dlygate4sd1_1 output227 (.A(net235),
    .X(branch_target_o[1]));
 sky130_fd_sc_hs__dlygate4sd1_1 output228 (.A(net236),
    .X(branch_target_o[20]));
 sky130_fd_sc_hs__dlygate4sd1_1 output229 (.A(net237),
    .X(branch_target_o[21]));
 sky130_fd_sc_hs__dlygate4sd1_1 output230 (.A(net238),
    .X(branch_target_o[22]));
 sky130_fd_sc_hs__dlygate4sd1_1 output231 (.A(net239),
    .X(branch_target_o[23]));
 sky130_fd_sc_hs__dlygate4sd1_1 output232 (.A(net240),
    .X(branch_target_o[24]));
 sky130_fd_sc_hs__dlygate4sd1_1 output233 (.A(net241),
    .X(branch_target_o[25]));
 sky130_fd_sc_hs__dlygate4sd1_1 output234 (.A(net242),
    .X(branch_target_o[26]));
 sky130_fd_sc_hs__dlygate4sd1_1 output235 (.A(net243),
    .X(branch_target_o[27]));
 sky130_fd_sc_hs__dlygate4sd1_1 output236 (.A(net244),
    .X(branch_target_o[28]));
 sky130_fd_sc_hs__dlygate4sd1_1 output237 (.A(net245),
    .X(branch_target_o[29]));
 sky130_fd_sc_hs__dlygate4sd1_1 output238 (.A(net246),
    .X(branch_target_o[2]));
 sky130_fd_sc_hs__dlygate4sd1_1 output239 (.A(net247),
    .X(branch_target_o[30]));
 sky130_fd_sc_hs__dlygate4sd1_1 output240 (.A(net248),
    .X(branch_target_o[31]));
 sky130_fd_sc_hs__dlygate4sd1_1 output241 (.A(net249),
    .X(branch_target_o[3]));
 sky130_fd_sc_hs__dlygate4sd1_1 output242 (.A(net250),
    .X(branch_target_o[4]));
 sky130_fd_sc_hs__dlygate4sd1_1 output243 (.A(net251),
    .X(branch_target_o[5]));
 sky130_fd_sc_hs__dlygate4sd1_1 output244 (.A(net252),
    .X(branch_target_o[6]));
 sky130_fd_sc_hs__dlygate4sd1_1 output245 (.A(net253),
    .X(branch_target_o[7]));
 sky130_fd_sc_hs__dlygate4sd1_1 output246 (.A(net254),
    .X(branch_target_o[8]));
 sky130_fd_sc_hs__dlygate4sd1_1 output247 (.A(net255),
    .X(branch_target_o[9]));
 sky130_fd_sc_hs__dlygate4sd1_1 output248 (.A(net256),
    .X(ex_valid_o));
 sky130_fd_sc_hs__dlygate4sd1_1 output249 (.A(net257),
    .X(imd_val_d_o[0]));
 sky130_fd_sc_hs__dlygate4sd1_1 output250 (.A(net258),
    .X(imd_val_d_o[10]));
 sky130_fd_sc_hs__dlygate4sd1_1 output251 (.A(net259),
    .X(imd_val_d_o[11]));
 sky130_fd_sc_hs__dlygate4sd1_1 output252 (.A(net260),
    .X(imd_val_d_o[12]));
 sky130_fd_sc_hs__dlygate4sd1_1 output253 (.A(net261),
    .X(imd_val_d_o[13]));
 sky130_fd_sc_hs__dlygate4sd1_1 output254 (.A(net262),
    .X(imd_val_d_o[14]));
 sky130_fd_sc_hs__dlygate4sd1_1 output255 (.A(net263),
    .X(imd_val_d_o[15]));
 sky130_fd_sc_hs__dlygate4sd1_1 output256 (.A(net264),
    .X(imd_val_d_o[16]));
 sky130_fd_sc_hs__dlygate4sd1_1 output257 (.A(net265),
    .X(imd_val_d_o[17]));
 sky130_fd_sc_hs__dlygate4sd1_1 output258 (.A(net266),
    .X(imd_val_d_o[18]));
 sky130_fd_sc_hs__dlygate4sd1_1 output259 (.A(net267),
    .X(imd_val_d_o[19]));
 sky130_fd_sc_hs__dlygate4sd1_1 output260 (.A(net268),
    .X(imd_val_d_o[1]));
 sky130_fd_sc_hs__dlygate4sd1_1 output261 (.A(net269),
    .X(imd_val_d_o[20]));
 sky130_fd_sc_hs__dlygate4sd1_1 output262 (.A(net270),
    .X(imd_val_d_o[21]));
 sky130_fd_sc_hs__dlygate4sd1_1 output263 (.A(net271),
    .X(imd_val_d_o[22]));
 sky130_fd_sc_hs__dlygate4sd1_1 output264 (.A(net272),
    .X(imd_val_d_o[23]));
 sky130_fd_sc_hs__dlygate4sd1_1 output265 (.A(net273),
    .X(imd_val_d_o[24]));
 sky130_fd_sc_hs__dlygate4sd1_1 output266 (.A(net274),
    .X(imd_val_d_o[25]));
 sky130_fd_sc_hs__dlygate4sd1_1 output267 (.A(net275),
    .X(imd_val_d_o[26]));
 sky130_fd_sc_hs__dlygate4sd1_1 output268 (.A(net276),
    .X(imd_val_d_o[27]));
 sky130_fd_sc_hs__dlygate4sd1_1 output269 (.A(net277),
    .X(imd_val_d_o[28]));
 sky130_fd_sc_hs__dlygate4sd1_1 output270 (.A(net278),
    .X(imd_val_d_o[29]));
 sky130_fd_sc_hs__dlygate4sd1_1 output271 (.A(net279),
    .X(imd_val_d_o[2]));
 sky130_fd_sc_hs__dlygate4sd1_1 output272 (.A(net280),
    .X(imd_val_d_o[30]));
 sky130_fd_sc_hs__dlygate4sd1_1 output273 (.A(net281),
    .X(imd_val_d_o[31]));
 sky130_fd_sc_hs__dlygate4sd1_1 output274 (.A(net282),
    .X(imd_val_d_o[34]));
 sky130_fd_sc_hs__dlygate4sd1_1 output275 (.A(net283),
    .X(imd_val_d_o[35]));
 sky130_fd_sc_hs__dlygate4sd1_1 output276 (.A(net284),
    .X(imd_val_d_o[36]));
 sky130_fd_sc_hs__dlygate4sd1_1 output277 (.A(net285),
    .X(imd_val_d_o[37]));
 sky130_fd_sc_hs__dlygate4sd1_1 output278 (.A(net286),
    .X(imd_val_d_o[38]));
 sky130_fd_sc_hs__dlygate4sd1_1 output279 (.A(net287),
    .X(imd_val_d_o[39]));
 sky130_fd_sc_hs__dlygate4sd1_1 output280 (.A(net288),
    .X(imd_val_d_o[3]));
 sky130_fd_sc_hs__dlygate4sd1_1 output281 (.A(net289),
    .X(imd_val_d_o[40]));
 sky130_fd_sc_hs__dlygate4sd1_1 output282 (.A(net290),
    .X(imd_val_d_o[41]));
 sky130_fd_sc_hs__dlygate4sd1_1 output283 (.A(net291),
    .X(imd_val_d_o[42]));
 sky130_fd_sc_hs__dlygate4sd1_1 output284 (.A(net292),
    .X(imd_val_d_o[43]));
 sky130_fd_sc_hs__dlygate4sd1_1 output285 (.A(net293),
    .X(imd_val_d_o[44]));
 sky130_fd_sc_hs__dlygate4sd1_1 output286 (.A(net294),
    .X(imd_val_d_o[45]));
 sky130_fd_sc_hs__dlygate4sd1_1 output287 (.A(net295),
    .X(imd_val_d_o[46]));
 sky130_fd_sc_hs__dlygate4sd1_1 output288 (.A(net296),
    .X(imd_val_d_o[47]));
 sky130_fd_sc_hs__dlygate4sd1_1 output289 (.A(net297),
    .X(imd_val_d_o[48]));
 sky130_fd_sc_hs__dlygate4sd1_1 output290 (.A(net298),
    .X(imd_val_d_o[49]));
 sky130_fd_sc_hs__dlygate4sd1_1 output291 (.A(net299),
    .X(imd_val_d_o[4]));
 sky130_fd_sc_hs__dlygate4sd1_1 output292 (.A(net300),
    .X(imd_val_d_o[50]));
 sky130_fd_sc_hs__dlygate4sd1_1 output293 (.A(net301),
    .X(imd_val_d_o[51]));
 sky130_fd_sc_hs__dlygate4sd1_1 output294 (.A(net302),
    .X(imd_val_d_o[52]));
 sky130_fd_sc_hs__dlygate4sd1_1 output295 (.A(net303),
    .X(imd_val_d_o[53]));
 sky130_fd_sc_hs__dlygate4sd1_1 output296 (.A(net304),
    .X(imd_val_d_o[54]));
 sky130_fd_sc_hs__dlygate4sd1_1 output297 (.A(net305),
    .X(imd_val_d_o[55]));
 sky130_fd_sc_hs__dlygate4sd1_1 output298 (.A(net306),
    .X(imd_val_d_o[56]));
 sky130_fd_sc_hs__dlygate4sd1_1 output299 (.A(net307),
    .X(imd_val_d_o[57]));
 sky130_fd_sc_hs__dlygate4sd1_1 output300 (.A(net308),
    .X(imd_val_d_o[58]));
 sky130_fd_sc_hs__dlygate4sd1_1 output301 (.A(net309),
    .X(imd_val_d_o[59]));
 sky130_fd_sc_hs__dlygate4sd1_1 output302 (.A(net310),
    .X(imd_val_d_o[5]));
 sky130_fd_sc_hs__dlygate4sd1_1 output303 (.A(net311),
    .X(imd_val_d_o[60]));
 sky130_fd_sc_hs__dlygate4sd1_1 output304 (.A(net312),
    .X(imd_val_d_o[61]));
 sky130_fd_sc_hs__dlygate4sd1_1 output305 (.A(net313),
    .X(imd_val_d_o[62]));
 sky130_fd_sc_hs__dlygate4sd1_1 output306 (.A(net314),
    .X(imd_val_d_o[63]));
 sky130_fd_sc_hs__dlygate4sd1_1 output307 (.A(net315),
    .X(imd_val_d_o[64]));
 sky130_fd_sc_hs__dlygate4sd1_1 output308 (.A(net316),
    .X(imd_val_d_o[65]));
 sky130_fd_sc_hs__dlygate4sd1_1 output309 (.A(net317),
    .X(imd_val_d_o[66]));
 sky130_fd_sc_hs__dlygate4sd1_1 output310 (.A(net318),
    .X(imd_val_d_o[67]));
 sky130_fd_sc_hs__dlygate4sd1_1 output311 (.A(net319),
    .X(imd_val_d_o[6]));
 sky130_fd_sc_hs__dlygate4sd1_1 output312 (.A(net320),
    .X(imd_val_d_o[7]));
 sky130_fd_sc_hs__dlygate4sd1_1 output313 (.A(net321),
    .X(imd_val_d_o[8]));
 sky130_fd_sc_hs__dlygate4sd1_1 output314 (.A(net322),
    .X(imd_val_d_o[9]));
 sky130_fd_sc_hs__dlygate4sd1_1 output315 (.A(net323),
    .X(imd_val_we_o[0]));
 sky130_fd_sc_hs__dlygate4sd1_1 output316 (.A(net324),
    .X(imd_val_we_o[1]));
 sky130_fd_sc_hs__dlygate4sd1_1 output317 (.A(net325),
    .X(result_ex_o[0]));
 sky130_fd_sc_hs__dlygate4sd1_1 output318 (.A(net326),
    .X(result_ex_o[10]));
 sky130_fd_sc_hs__dlygate4sd1_1 output319 (.A(net327),
    .X(result_ex_o[11]));
 sky130_fd_sc_hs__dlygate4sd1_1 output320 (.A(net328),
    .X(result_ex_o[12]));
 sky130_fd_sc_hs__dlygate4sd1_1 output321 (.A(net329),
    .X(result_ex_o[13]));
 sky130_fd_sc_hs__dlygate4sd1_1 output322 (.A(net330),
    .X(result_ex_o[14]));
 sky130_fd_sc_hs__dlygate4sd1_1 output323 (.A(net331),
    .X(result_ex_o[15]));
 sky130_fd_sc_hs__dlygate4sd1_1 output324 (.A(net332),
    .X(result_ex_o[16]));
 sky130_fd_sc_hs__dlygate4sd1_1 output325 (.A(net333),
    .X(result_ex_o[17]));
 sky130_fd_sc_hs__dlygate4sd1_1 output326 (.A(net334),
    .X(result_ex_o[18]));
 sky130_fd_sc_hs__dlygate4sd1_1 output327 (.A(net335),
    .X(result_ex_o[19]));
 sky130_fd_sc_hs__dlygate4sd1_1 output328 (.A(net336),
    .X(result_ex_o[1]));
 sky130_fd_sc_hs__dlygate4sd1_1 output329 (.A(net337),
    .X(result_ex_o[20]));
 sky130_fd_sc_hs__dlygate4sd1_1 output330 (.A(net338),
    .X(result_ex_o[21]));
 sky130_fd_sc_hs__dlygate4sd1_1 output331 (.A(net339),
    .X(result_ex_o[22]));
 sky130_fd_sc_hs__dlygate4sd1_1 output332 (.A(net340),
    .X(result_ex_o[23]));
 sky130_fd_sc_hs__dlygate4sd1_1 output333 (.A(net341),
    .X(result_ex_o[24]));
 sky130_fd_sc_hs__dlygate4sd1_1 output334 (.A(net342),
    .X(result_ex_o[25]));
 sky130_fd_sc_hs__dlygate4sd1_1 output335 (.A(net343),
    .X(result_ex_o[26]));
 sky130_fd_sc_hs__dlygate4sd1_1 output336 (.A(net344),
    .X(result_ex_o[27]));
 sky130_fd_sc_hs__dlygate4sd1_1 output337 (.A(net345),
    .X(result_ex_o[28]));
 sky130_fd_sc_hs__dlygate4sd1_1 output338 (.A(net346),
    .X(result_ex_o[29]));
 sky130_fd_sc_hs__dlygate4sd1_1 output339 (.A(net347),
    .X(result_ex_o[2]));
 sky130_fd_sc_hs__dlygate4sd1_1 output340 (.A(net348),
    .X(result_ex_o[30]));
 sky130_fd_sc_hs__dlygate4sd1_1 output341 (.A(net349),
    .X(result_ex_o[31]));
 sky130_fd_sc_hs__dlygate4sd1_1 output342 (.A(net350),
    .X(result_ex_o[3]));
 sky130_fd_sc_hs__dlygate4sd1_1 output343 (.A(net351),
    .X(result_ex_o[4]));
 sky130_fd_sc_hs__dlygate4sd1_1 output344 (.A(net352),
    .X(result_ex_o[5]));
 sky130_fd_sc_hs__dlygate4sd1_1 output345 (.A(net353),
    .X(result_ex_o[6]));
 sky130_fd_sc_hs__dlygate4sd1_1 output346 (.A(net354),
    .X(result_ex_o[7]));
 sky130_fd_sc_hs__dlygate4sd1_1 output347 (.A(net355),
    .X(result_ex_o[8]));
 sky130_fd_sc_hs__dlygate4sd1_1 output348 (.A(net356),
    .X(result_ex_o[9]));
 sky130_fd_sc_hs__dlygate4sd1_1 max_cap349 (.A(net358),
    .X(net357));
 sky130_fd_sc_hs__dlygate4sd1_1 load_slew350 (.A(net359),
    .X(net358));
 sky130_fd_sc_hs__dlygate4sd1_1 load_slew351 (.A(net360),
    .X(net359));
 sky130_fd_sc_hs__dlygate4sd1_1 load_slew352 (.A(net361),
    .X(net360));
 sky130_fd_sc_hs__dlygate4sd1_1 load_slew353 (.A(net362),
    .X(net361));
 sky130_fd_sc_hs__dlygate4sd1_1 load_slew354 (.A(net190),
    .X(net362));
 sky130_fd_sc_hs__conb_1 _7887__355 (.LO(net363));
 sky130_fd_sc_hs__conb_1 _7888__356 (.LO(net364));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_3_0_0_clk_i (.A(clknet_0_clk_i),
    .X(clknet_3_0_0_clk_i));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_3_1_0_clk_i (.A(clknet_0_clk_i),
    .X(clknet_3_1_0_clk_i));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_3_2_0_clk_i (.A(clknet_0_clk_i),
    .X(clknet_3_2_0_clk_i));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_3_3_0_clk_i (.A(clknet_0_clk_i),
    .X(clknet_3_3_0_clk_i));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_3_4_0_clk_i (.A(clknet_0_clk_i),
    .X(clknet_3_4_0_clk_i));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_3_5_0_clk_i (.A(clknet_0_clk_i),
    .X(clknet_3_5_0_clk_i));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_3_6_0_clk_i (.A(clknet_0_clk_i),
    .X(clknet_3_6_0_clk_i));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_3_7_0_clk_i (.A(clknet_0_clk_i),
    .X(clknet_3_7_0_clk_i));
 sky130_fd_sc_hs__clkinv_2 clkload0 (.A(clknet_3_1_0_clk_i));
 sky130_fd_sc_hs__clkinv_2 clkload1 (.A(clknet_3_2_0_clk_i));
 sky130_fd_sc_hs__clkinv_4 clkload2 (.A(clknet_3_3_0_clk_i));
 sky130_fd_sc_hs__inv_8 clkload3 (.A(clknet_3_4_0_clk_i));
 sky130_fd_sc_hs__clkinv_4 clkload4 (.A(clknet_3_5_0_clk_i));
 sky130_fd_sc_hs__inv_8 clkload5 (.A(clknet_3_6_0_clk_i));
 sky130_fd_sc_hs__clkinv_4 clkload6 (.A(clknet_3_7_0_clk_i));
 sky130_fd_sc_hs__buf_16 load_slew1 (.A(net193),
    .X(net365));
 sky130_fd_sc_hs__clkbuf_8 load_slew2 (.A(_0379_),
    .X(net366));
 sky130_fd_sc_hs__diode_2 ANTENNA_1 (.DIODE(net242));
 sky130_fd_sc_hs__diode_2 ANTENNA_2 (.DIODE(net242));
 sky130_fd_sc_hs__diode_2 ANTENNA_3 (.DIODE(net242));
 sky130_fd_sc_hs__diode_2 ANTENNA_4 (.DIODE(net242));
 sky130_fd_sc_hs__diode_2 ANTENNA_5 (.DIODE(net242));
 sky130_fd_sc_hs__diode_2 ANTENNA_6 (.DIODE(net242));
 sky130_fd_sc_hs__diode_2 ANTENNA_7 (.DIODE(net242));
 sky130_fd_sc_hs__diode_2 ANTENNA_8 (.DIODE(net243));
 sky130_fd_sc_hs__diode_2 ANTENNA_9 (.DIODE(net243));
 sky130_fd_sc_hs__diode_2 ANTENNA_10 (.DIODE(net245));
 sky130_fd_sc_hs__diode_2 ANTENNA_11 (.DIODE(net245));
 sky130_fd_sc_hs__diode_2 ANTENNA_12 (.DIODE(net245));
 sky130_fd_sc_hs__diode_2 ANTENNA_13 (.DIODE(net250));
 sky130_fd_sc_hs__diode_2 ANTENNA_14 (.DIODE(net250));
 sky130_fd_sc_hs__diode_2 ANTENNA_15 (.DIODE(net250));
 sky130_fd_sc_hs__diode_2 ANTENNA_16 (.DIODE(net250));
 sky130_fd_sc_hs__diode_2 ANTENNA_17 (.DIODE(net250));
 sky130_fd_sc_hs__diode_2 ANTENNA_18 (.DIODE(net250));
 sky130_fd_sc_hs__diode_2 ANTENNA_19 (.DIODE(net250));
 sky130_fd_sc_hs__diode_2 ANTENNA_20 (.DIODE(net310));
 sky130_fd_sc_hs__diode_2 ANTENNA_21 (.DIODE(imd_val_q_i[47]));
 sky130_fd_sc_hs__diode_2 ANTENNA_22 (.DIODE(net310));
 sky130_fd_sc_hs__diode_2 ANTENNA_23 (.DIODE(net310));
 sky130_fd_sc_hs__diode_2 ANTENNA_24 (.DIODE(net310));
 sky130_fd_sc_hs__diode_2 ANTENNA_25 (.DIODE(net310));
 sky130_fd_sc_hs__diode_2 ANTENNA_26 (.DIODE(net215));
 sky130_fd_sc_hs__diode_2 ANTENNA_27 (.DIODE(net266));
 sky130_fd_sc_hs__diode_2 ANTENNA_28 (.DIODE(net215));
 sky130_fd_sc_hs__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_0_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_46 ();
 sky130_fd_sc_hs__fill_4 FILLER_0_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_75 ();
 sky130_fd_sc_hs__fill_4 FILLER_0_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_104 ();
 sky130_fd_sc_hs__fill_4 FILLER_0_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_133 ();
 sky130_fd_sc_hs__fill_4 FILLER_0_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_162 ();
 sky130_fd_sc_hs__fill_4 FILLER_0_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_191 ();
 sky130_fd_sc_hs__fill_4 FILLER_0_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_220 ();
 sky130_fd_sc_hs__fill_4 FILLER_0_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_249 ();
 sky130_fd_sc_hs__fill_4 FILLER_0_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_278 ();
 sky130_fd_sc_hs__fill_4 FILLER_0_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_307 ();
 sky130_fd_sc_hs__fill_4 FILLER_0_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_336 ();
 sky130_fd_sc_hs__fill_4 FILLER_0_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_365 ();
 sky130_fd_sc_hs__fill_4 FILLER_0_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_394 ();
 sky130_fd_sc_hs__fill_4 FILLER_0_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_423 ();
 sky130_fd_sc_hs__fill_4 FILLER_0_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_452 ();
 sky130_fd_sc_hs__fill_4 FILLER_0_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_481 ();
 sky130_fd_sc_hs__fill_4 FILLER_0_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_510 ();
 sky130_fd_sc_hs__fill_4 FILLER_0_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_0_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_0_539 ();
 sky130_fd_sc_hs__fill_1 FILLER_1_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_9 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_17 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_25 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_33 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_41 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_49 ();
 sky130_fd_sc_hs__fill_1 FILLER_1_57 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_1_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_1_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_1_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_1_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_1_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_1_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_1_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_1_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_1_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_1_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_2_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_2_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_2_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_2_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_2_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_2_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_302 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_310 ();
 sky130_fd_sc_hs__fill_1 FILLER_2_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_2_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_2_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_2_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_2_526 ();
 sky130_fd_sc_hs__fill_4 FILLER_2_534 ();
 sky130_fd_sc_hs__fill_2 FILLER_2_538 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_3_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_3_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_3_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_3_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_3_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_3_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_3_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_3_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_3_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_3_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_3_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_4_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_4_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_4_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_4_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_4_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_4_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_302 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_310 ();
 sky130_fd_sc_hs__fill_1 FILLER_4_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_4_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_4_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_4_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_4_526 ();
 sky130_fd_sc_hs__fill_4 FILLER_4_534 ();
 sky130_fd_sc_hs__fill_2 FILLER_4_538 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_16 ();
 sky130_fd_sc_hs__fill_1 FILLER_5_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_27 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_35 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_43 ();
 sky130_fd_sc_hs__fill_4 FILLER_5_51 ();
 sky130_fd_sc_hs__fill_2 FILLER_5_55 ();
 sky130_fd_sc_hs__fill_1 FILLER_5_57 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_5_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_5_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_5_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_5_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_5_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_5_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_5_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_5_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_5_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_5_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_16 ();
 sky130_fd_sc_hs__fill_1 FILLER_6_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_6_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_6_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_6_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_6_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_302 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_310 ();
 sky130_fd_sc_hs__fill_1 FILLER_6_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_6_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_6_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_6_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_6_526 ();
 sky130_fd_sc_hs__fill_4 FILLER_6_534 ();
 sky130_fd_sc_hs__fill_2 FILLER_6_538 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_16 ();
 sky130_fd_sc_hs__fill_1 FILLER_7_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_33 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_41 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_49 ();
 sky130_fd_sc_hs__fill_1 FILLER_7_57 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_7_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_7_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_7_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_7_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_7_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_7_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_7_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_7_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_7_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_7_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_16 ();
 sky130_fd_sc_hs__fill_1 FILLER_8_24 ();
 sky130_fd_sc_hs__fill_2 FILLER_8_27 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_8_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_8_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_8_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_8_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_302 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_310 ();
 sky130_fd_sc_hs__fill_1 FILLER_8_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_8_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_8_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_8_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_8_526 ();
 sky130_fd_sc_hs__fill_4 FILLER_8_534 ();
 sky130_fd_sc_hs__fill_2 FILLER_8_538 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_16 ();
 sky130_fd_sc_hs__fill_1 FILLER_9_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_27 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_35 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_43 ();
 sky130_fd_sc_hs__fill_4 FILLER_9_51 ();
 sky130_fd_sc_hs__fill_2 FILLER_9_55 ();
 sky130_fd_sc_hs__fill_1 FILLER_9_57 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_9_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_9_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_9_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_9_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_9_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_9_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_9_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_9_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_9_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_9_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_10_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_10_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_10_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_10_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_10_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_10_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_302 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_310 ();
 sky130_fd_sc_hs__fill_1 FILLER_10_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_10_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_10_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_10_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_10_526 ();
 sky130_fd_sc_hs__fill_4 FILLER_10_534 ();
 sky130_fd_sc_hs__fill_2 FILLER_10_538 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_0 ();
 sky130_fd_sc_hs__fill_4 FILLER_11_8 ();
 sky130_fd_sc_hs__fill_2 FILLER_11_12 ();
 sky130_fd_sc_hs__fill_1 FILLER_11_14 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_23 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_31 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_39 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_47 ();
 sky130_fd_sc_hs__fill_2 FILLER_11_55 ();
 sky130_fd_sc_hs__fill_1 FILLER_11_57 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_11_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_11_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_191 ();
 sky130_fd_sc_hs__fill_1 FILLER_11_199 ();
 sky130_fd_sc_hs__fill_4 FILLER_11_203 ();
 sky130_fd_sc_hs__fill_2 FILLER_11_207 ();
 sky130_fd_sc_hs__fill_1 FILLER_11_209 ();
 sky130_fd_sc_hs__fill_1 FILLER_11_231 ();
 sky130_fd_sc_hs__fill_4 FILLER_11_236 ();
 sky130_fd_sc_hs__fill_1 FILLER_11_243 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_11_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_11_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_11_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_11_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_11_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_11_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_11_539 ();
 sky130_fd_sc_hs__fill_4 FILLER_12_0 ();
 sky130_fd_sc_hs__fill_1 FILLER_12_4 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_21 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_12_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_12_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_170 ();
 sky130_fd_sc_hs__fill_4 FILLER_12_178 ();
 sky130_fd_sc_hs__fill_2 FILLER_12_182 ();
 sky130_fd_sc_hs__fill_1 FILLER_12_202 ();
 sky130_fd_sc_hs__fill_2 FILLER_12_259 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_275 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_283 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_307 ();
 sky130_fd_sc_hs__fill_4 FILLER_12_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_12_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_12_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_12_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_12_526 ();
 sky130_fd_sc_hs__fill_4 FILLER_12_534 ();
 sky130_fd_sc_hs__fill_2 FILLER_12_538 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_13_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_13_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_13_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_175 ();
 sky130_fd_sc_hs__fill_4 FILLER_13_183 ();
 sky130_fd_sc_hs__fill_1 FILLER_13_187 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_194 ();
 sky130_fd_sc_hs__fill_2 FILLER_13_230 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_241 ();
 sky130_fd_sc_hs__fill_2 FILLER_13_267 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_13_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_13_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_13_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_13_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_13_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_13_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_14_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_14_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_14_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_14_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_162 ();
 sky130_fd_sc_hs__fill_2 FILLER_14_170 ();
 sky130_fd_sc_hs__fill_1 FILLER_14_204 ();
 sky130_fd_sc_hs__fill_1 FILLER_14_208 ();
 sky130_fd_sc_hs__fill_1 FILLER_14_248 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_14_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_262 ();
 sky130_fd_sc_hs__fill_2 FILLER_14_297 ();
 sky130_fd_sc_hs__fill_1 FILLER_14_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_305 ();
 sky130_fd_sc_hs__fill_4 FILLER_14_313 ();
 sky130_fd_sc_hs__fill_2 FILLER_14_317 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_14_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_14_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_14_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_14_526 ();
 sky130_fd_sc_hs__fill_4 FILLER_14_534 ();
 sky130_fd_sc_hs__fill_2 FILLER_14_538 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_0 ();
 sky130_fd_sc_hs__fill_2 FILLER_15_8 ();
 sky130_fd_sc_hs__fill_1 FILLER_15_10 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_19 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_27 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_35 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_43 ();
 sky130_fd_sc_hs__fill_4 FILLER_15_51 ();
 sky130_fd_sc_hs__fill_2 FILLER_15_55 ();
 sky130_fd_sc_hs__fill_1 FILLER_15_57 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_15_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_141 ();
 sky130_fd_sc_hs__fill_2 FILLER_15_149 ();
 sky130_fd_sc_hs__fill_1 FILLER_15_154 ();
 sky130_fd_sc_hs__fill_1 FILLER_15_173 ();
 sky130_fd_sc_hs__fill_2 FILLER_15_175 ();
 sky130_fd_sc_hs__fill_2 FILLER_15_180 ();
 sky130_fd_sc_hs__fill_1 FILLER_15_182 ();
 sky130_fd_sc_hs__fill_2 FILLER_15_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_196 ();
 sky130_fd_sc_hs__fill_2 FILLER_15_204 ();
 sky130_fd_sc_hs__fill_1 FILLER_15_206 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_220 ();
 sky130_fd_sc_hs__fill_4 FILLER_15_228 ();
 sky130_fd_sc_hs__fill_2 FILLER_15_238 ();
 sky130_fd_sc_hs__fill_1 FILLER_15_240 ();
 sky130_fd_sc_hs__fill_4 FILLER_15_245 ();
 sky130_fd_sc_hs__fill_1 FILLER_15_249 ();
 sky130_fd_sc_hs__fill_1 FILLER_15_253 ();
 sky130_fd_sc_hs__fill_4 FILLER_15_257 ();
 sky130_fd_sc_hs__fill_2 FILLER_15_261 ();
 sky130_fd_sc_hs__fill_4 FILLER_15_267 ();
 sky130_fd_sc_hs__fill_2 FILLER_15_282 ();
 sky130_fd_sc_hs__fill_1 FILLER_15_284 ();
 sky130_fd_sc_hs__fill_2 FILLER_15_288 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_312 ();
 sky130_fd_sc_hs__fill_4 FILLER_15_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_329 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_337 ();
 sky130_fd_sc_hs__fill_2 FILLER_15_345 ();
 sky130_fd_sc_hs__fill_1 FILLER_15_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_15_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_15_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_15_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_15_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_15_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_16_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_16_28 ();
 sky130_fd_sc_hs__fill_1 FILLER_16_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_39 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_47 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_55 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_63 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_71 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_79 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_16_144 ();
 sky130_fd_sc_hs__fill_2 FILLER_16_164 ();
 sky130_fd_sc_hs__fill_1 FILLER_16_166 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_170 ();
 sky130_fd_sc_hs__fill_2 FILLER_16_178 ();
 sky130_fd_sc_hs__fill_4 FILLER_16_183 ();
 sky130_fd_sc_hs__fill_2 FILLER_16_187 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_192 ();
 sky130_fd_sc_hs__fill_2 FILLER_16_200 ();
 sky130_fd_sc_hs__fill_1 FILLER_16_202 ();
 sky130_fd_sc_hs__fill_4 FILLER_16_204 ();
 sky130_fd_sc_hs__fill_4 FILLER_16_211 ();
 sky130_fd_sc_hs__fill_1 FILLER_16_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_219 ();
 sky130_fd_sc_hs__fill_4 FILLER_16_227 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_234 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_242 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_250 ();
 sky130_fd_sc_hs__fill_2 FILLER_16_258 ();
 sky130_fd_sc_hs__fill_1 FILLER_16_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_278 ();
 sky130_fd_sc_hs__fill_4 FILLER_16_286 ();
 sky130_fd_sc_hs__fill_1 FILLER_16_290 ();
 sky130_fd_sc_hs__fill_2 FILLER_16_294 ();
 sky130_fd_sc_hs__fill_1 FILLER_16_296 ();
 sky130_fd_sc_hs__fill_4 FILLER_16_300 ();
 sky130_fd_sc_hs__fill_2 FILLER_16_304 ();
 sky130_fd_sc_hs__fill_1 FILLER_16_306 ();
 sky130_fd_sc_hs__fill_2 FILLER_16_310 ();
 sky130_fd_sc_hs__fill_4 FILLER_16_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_341 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_365 ();
 sky130_fd_sc_hs__fill_4 FILLER_16_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_16_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_16_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_16_526 ();
 sky130_fd_sc_hs__fill_4 FILLER_16_534 ();
 sky130_fd_sc_hs__fill_2 FILLER_16_538 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_0 ();
 sky130_fd_sc_hs__fill_4 FILLER_17_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_20 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_36 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_44 ();
 sky130_fd_sc_hs__fill_4 FILLER_17_52 ();
 sky130_fd_sc_hs__fill_2 FILLER_17_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_17_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_141 ();
 sky130_fd_sc_hs__fill_1 FILLER_17_149 ();
 sky130_fd_sc_hs__fill_1 FILLER_17_156 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_163 ();
 sky130_fd_sc_hs__fill_2 FILLER_17_171 ();
 sky130_fd_sc_hs__fill_1 FILLER_17_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_193 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_222 ();
 sky130_fd_sc_hs__fill_2 FILLER_17_230 ();
 sky130_fd_sc_hs__fill_2 FILLER_17_242 ();
 sky130_fd_sc_hs__fill_1 FILLER_17_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_272 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_280 ();
 sky130_fd_sc_hs__fill_2 FILLER_17_288 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_317 ();
 sky130_fd_sc_hs__fill_4 FILLER_17_328 ();
 sky130_fd_sc_hs__fill_2 FILLER_17_337 ();
 sky130_fd_sc_hs__fill_1 FILLER_17_339 ();
 sky130_fd_sc_hs__fill_4 FILLER_17_343 ();
 sky130_fd_sc_hs__fill_1 FILLER_17_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_17_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_17_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_17_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_17_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_17_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_18_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_18_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_18_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_18_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_146 ();
 sky130_fd_sc_hs__fill_2 FILLER_18_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_166 ();
 sky130_fd_sc_hs__fill_2 FILLER_18_174 ();
 sky130_fd_sc_hs__fill_1 FILLER_18_176 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_180 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_188 ();
 sky130_fd_sc_hs__fill_4 FILLER_18_196 ();
 sky130_fd_sc_hs__fill_2 FILLER_18_200 ();
 sky130_fd_sc_hs__fill_1 FILLER_18_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_220 ();
 sky130_fd_sc_hs__fill_2 FILLER_18_228 ();
 sky130_fd_sc_hs__fill_1 FILLER_18_230 ();
 sky130_fd_sc_hs__fill_4 FILLER_18_249 ();
 sky130_fd_sc_hs__fill_2 FILLER_18_253 ();
 sky130_fd_sc_hs__fill_2 FILLER_18_258 ();
 sky130_fd_sc_hs__fill_1 FILLER_18_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_286 ();
 sky130_fd_sc_hs__fill_4 FILLER_18_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_301 ();
 sky130_fd_sc_hs__fill_4 FILLER_18_309 ();
 sky130_fd_sc_hs__fill_2 FILLER_18_316 ();
 sky130_fd_sc_hs__fill_1 FILLER_18_318 ();
 sky130_fd_sc_hs__fill_1 FILLER_18_320 ();
 sky130_fd_sc_hs__fill_4 FILLER_18_345 ();
 sky130_fd_sc_hs__fill_2 FILLER_18_349 ();
 sky130_fd_sc_hs__fill_1 FILLER_18_351 ();
 sky130_fd_sc_hs__fill_4 FILLER_18_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_364 ();
 sky130_fd_sc_hs__fill_4 FILLER_18_372 ();
 sky130_fd_sc_hs__fill_1 FILLER_18_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_18_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_18_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_18_526 ();
 sky130_fd_sc_hs__fill_4 FILLER_18_534 ();
 sky130_fd_sc_hs__fill_2 FILLER_18_538 ();
 sky130_fd_sc_hs__fill_1 FILLER_19_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_17 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_25 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_33 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_41 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_49 ();
 sky130_fd_sc_hs__fill_1 FILLER_19_57 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_19_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_125 ();
 sky130_fd_sc_hs__fill_1 FILLER_19_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_137 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_145 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_153 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_161 ();
 sky130_fd_sc_hs__fill_4 FILLER_19_169 ();
 sky130_fd_sc_hs__fill_1 FILLER_19_173 ();
 sky130_fd_sc_hs__fill_4 FILLER_19_175 ();
 sky130_fd_sc_hs__fill_1 FILLER_19_179 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_191 ();
 sky130_fd_sc_hs__fill_4 FILLER_19_199 ();
 sky130_fd_sc_hs__fill_1 FILLER_19_203 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_19_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_233 ();
 sky130_fd_sc_hs__fill_4 FILLER_19_241 ();
 sky130_fd_sc_hs__fill_2 FILLER_19_245 ();
 sky130_fd_sc_hs__fill_1 FILLER_19_247 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_251 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_259 ();
 sky130_fd_sc_hs__fill_4 FILLER_19_267 ();
 sky130_fd_sc_hs__fill_1 FILLER_19_271 ();
 sky130_fd_sc_hs__fill_4 FILLER_19_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_305 ();
 sky130_fd_sc_hs__fill_1 FILLER_19_313 ();
 sky130_fd_sc_hs__fill_1 FILLER_19_332 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_336 ();
 sky130_fd_sc_hs__fill_1 FILLER_19_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_367 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_375 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_383 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_391 ();
 sky130_fd_sc_hs__fill_4 FILLER_19_399 ();
 sky130_fd_sc_hs__fill_2 FILLER_19_403 ();
 sky130_fd_sc_hs__fill_1 FILLER_19_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_19_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_19_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_19_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_19_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_20_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_20_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_20_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_120 ();
 sky130_fd_sc_hs__fill_4 FILLER_20_128 ();
 sky130_fd_sc_hs__fill_1 FILLER_20_138 ();
 sky130_fd_sc_hs__fill_1 FILLER_20_144 ();
 sky130_fd_sc_hs__fill_4 FILLER_20_146 ();
 sky130_fd_sc_hs__fill_2 FILLER_20_150 ();
 sky130_fd_sc_hs__fill_1 FILLER_20_152 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_156 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_164 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_172 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_180 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_188 ();
 sky130_fd_sc_hs__fill_4 FILLER_20_196 ();
 sky130_fd_sc_hs__fill_2 FILLER_20_200 ();
 sky130_fd_sc_hs__fill_1 FILLER_20_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_220 ();
 sky130_fd_sc_hs__fill_2 FILLER_20_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_249 ();
 sky130_fd_sc_hs__fill_4 FILLER_20_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_262 ();
 sky130_fd_sc_hs__fill_2 FILLER_20_270 ();
 sky130_fd_sc_hs__fill_1 FILLER_20_272 ();
 sky130_fd_sc_hs__fill_4 FILLER_20_280 ();
 sky130_fd_sc_hs__fill_2 FILLER_20_284 ();
 sky130_fd_sc_hs__fill_1 FILLER_20_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_293 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_301 ();
 sky130_fd_sc_hs__fill_2 FILLER_20_309 ();
 sky130_fd_sc_hs__fill_1 FILLER_20_311 ();
 sky130_fd_sc_hs__fill_1 FILLER_20_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_320 ();
 sky130_fd_sc_hs__fill_2 FILLER_20_328 ();
 sky130_fd_sc_hs__fill_1 FILLER_20_330 ();
 sky130_fd_sc_hs__fill_4 FILLER_20_334 ();
 sky130_fd_sc_hs__fill_1 FILLER_20_338 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_20_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_20_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_20_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_20_526 ();
 sky130_fd_sc_hs__fill_4 FILLER_20_534 ();
 sky130_fd_sc_hs__fill_2 FILLER_20_538 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_21_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_21_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_117 ();
 sky130_fd_sc_hs__fill_1 FILLER_21_125 ();
 sky130_fd_sc_hs__fill_1 FILLER_21_144 ();
 sky130_fd_sc_hs__fill_4 FILLER_21_166 ();
 sky130_fd_sc_hs__fill_1 FILLER_21_170 ();
 sky130_fd_sc_hs__fill_4 FILLER_21_193 ();
 sky130_fd_sc_hs__fill_2 FILLER_21_197 ();
 sky130_fd_sc_hs__fill_1 FILLER_21_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_219 ();
 sky130_fd_sc_hs__fill_4 FILLER_21_227 ();
 sky130_fd_sc_hs__fill_1 FILLER_21_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_265 ();
 sky130_fd_sc_hs__fill_1 FILLER_21_273 ();
 sky130_fd_sc_hs__fill_1 FILLER_21_277 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_21_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_299 ();
 sky130_fd_sc_hs__fill_2 FILLER_21_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_319 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_327 ();
 sky130_fd_sc_hs__fill_2 FILLER_21_335 ();
 sky130_fd_sc_hs__fill_2 FILLER_21_346 ();
 sky130_fd_sc_hs__fill_4 FILLER_21_349 ();
 sky130_fd_sc_hs__fill_2 FILLER_21_353 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_358 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_366 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_374 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_382 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_390 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_398 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_21_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_21_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_21_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_21_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_22_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_22_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_22_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_112 ();
 sky130_fd_sc_hs__fill_2 FILLER_22_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_130 ();
 sky130_fd_sc_hs__fill_4 FILLER_22_138 ();
 sky130_fd_sc_hs__fill_2 FILLER_22_142 ();
 sky130_fd_sc_hs__fill_1 FILLER_22_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_164 ();
 sky130_fd_sc_hs__fill_4 FILLER_22_172 ();
 sky130_fd_sc_hs__fill_1 FILLER_22_176 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_180 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_188 ();
 sky130_fd_sc_hs__fill_1 FILLER_22_196 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_243 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_251 ();
 sky130_fd_sc_hs__fill_2 FILLER_22_259 ();
 sky130_fd_sc_hs__fill_2 FILLER_22_262 ();
 sky130_fd_sc_hs__fill_1 FILLER_22_264 ();
 sky130_fd_sc_hs__fill_1 FILLER_22_268 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_287 ();
 sky130_fd_sc_hs__fill_1 FILLER_22_295 ();
 sky130_fd_sc_hs__fill_1 FILLER_22_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_320 ();
 sky130_fd_sc_hs__fill_4 FILLER_22_328 ();
 sky130_fd_sc_hs__fill_1 FILLER_22_332 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_343 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_351 ();
 sky130_fd_sc_hs__fill_4 FILLER_22_359 ();
 sky130_fd_sc_hs__fill_2 FILLER_22_363 ();
 sky130_fd_sc_hs__fill_1 FILLER_22_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_369 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_22_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_22_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_22_526 ();
 sky130_fd_sc_hs__fill_4 FILLER_22_534 ();
 sky130_fd_sc_hs__fill_2 FILLER_22_538 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_8 ();
 sky130_fd_sc_hs__fill_4 FILLER_23_16 ();
 sky130_fd_sc_hs__fill_2 FILLER_23_20 ();
 sky130_fd_sc_hs__fill_1 FILLER_23_22 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_31 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_39 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_47 ();
 sky130_fd_sc_hs__fill_2 FILLER_23_55 ();
 sky130_fd_sc_hs__fill_1 FILLER_23_57 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_99 ();
 sky130_fd_sc_hs__fill_2 FILLER_23_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_23_109 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_135 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_143 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_164 ();
 sky130_fd_sc_hs__fill_2 FILLER_23_172 ();
 sky130_fd_sc_hs__fill_1 FILLER_23_175 ();
 sky130_fd_sc_hs__fill_2 FILLER_23_194 ();
 sky130_fd_sc_hs__fill_4 FILLER_23_236 ();
 sky130_fd_sc_hs__fill_2 FILLER_23_240 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_261 ();
 sky130_fd_sc_hs__fill_1 FILLER_23_269 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_23_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_302 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_310 ();
 sky130_fd_sc_hs__fill_2 FILLER_23_318 ();
 sky130_fd_sc_hs__fill_1 FILLER_23_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_23_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_357 ();
 sky130_fd_sc_hs__fill_2 FILLER_23_365 ();
 sky130_fd_sc_hs__fill_1 FILLER_23_367 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_394 ();
 sky130_fd_sc_hs__fill_4 FILLER_23_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_23_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_23_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_23_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_23_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_8 ();
 sky130_fd_sc_hs__fill_4 FILLER_24_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_24_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_70 ();
 sky130_fd_sc_hs__fill_2 FILLER_24_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_24_80 ();
 sky130_fd_sc_hs__fill_2 FILLER_24_84 ();
 sky130_fd_sc_hs__fill_1 FILLER_24_86 ();
 sky130_fd_sc_hs__fill_1 FILLER_24_88 ();
 sky130_fd_sc_hs__fill_4 FILLER_24_107 ();
 sky130_fd_sc_hs__fill_2 FILLER_24_111 ();
 sky130_fd_sc_hs__fill_1 FILLER_24_113 ();
 sky130_fd_sc_hs__fill_4 FILLER_24_117 ();
 sky130_fd_sc_hs__fill_2 FILLER_24_121 ();
 sky130_fd_sc_hs__fill_1 FILLER_24_144 ();
 sky130_fd_sc_hs__fill_4 FILLER_24_146 ();
 sky130_fd_sc_hs__fill_1 FILLER_24_150 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_154 ();
 sky130_fd_sc_hs__fill_2 FILLER_24_162 ();
 sky130_fd_sc_hs__fill_1 FILLER_24_164 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_168 ();
 sky130_fd_sc_hs__fill_4 FILLER_24_176 ();
 sky130_fd_sc_hs__fill_2 FILLER_24_180 ();
 sky130_fd_sc_hs__fill_4 FILLER_24_185 ();
 sky130_fd_sc_hs__fill_1 FILLER_24_189 ();
 sky130_fd_sc_hs__fill_4 FILLER_24_193 ();
 sky130_fd_sc_hs__fill_2 FILLER_24_214 ();
 sky130_fd_sc_hs__fill_1 FILLER_24_216 ();
 sky130_fd_sc_hs__fill_1 FILLER_24_238 ();
 sky130_fd_sc_hs__fill_1 FILLER_24_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_270 ();
 sky130_fd_sc_hs__fill_2 FILLER_24_283 ();
 sky130_fd_sc_hs__fill_1 FILLER_24_285 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_307 ();
 sky130_fd_sc_hs__fill_4 FILLER_24_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_344 ();
 sky130_fd_sc_hs__fill_1 FILLER_24_352 ();
 sky130_fd_sc_hs__fill_4 FILLER_24_366 ();
 sky130_fd_sc_hs__fill_2 FILLER_24_370 ();
 sky130_fd_sc_hs__fill_4 FILLER_24_378 ();
 sky130_fd_sc_hs__fill_1 FILLER_24_382 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_24_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_24_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_24_526 ();
 sky130_fd_sc_hs__fill_4 FILLER_24_534 ();
 sky130_fd_sc_hs__fill_2 FILLER_24_538 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_25_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_83 ();
 sky130_fd_sc_hs__fill_4 FILLER_25_91 ();
 sky130_fd_sc_hs__fill_1 FILLER_25_95 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_101 ();
 sky130_fd_sc_hs__fill_4 FILLER_25_109 ();
 sky130_fd_sc_hs__fill_2 FILLER_25_113 ();
 sky130_fd_sc_hs__fill_1 FILLER_25_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_128 ();
 sky130_fd_sc_hs__fill_1 FILLER_25_136 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_156 ();
 sky130_fd_sc_hs__fill_4 FILLER_25_164 ();
 sky130_fd_sc_hs__fill_2 FILLER_25_168 ();
 sky130_fd_sc_hs__fill_1 FILLER_25_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_175 ();
 sky130_fd_sc_hs__fill_4 FILLER_25_183 ();
 sky130_fd_sc_hs__fill_1 FILLER_25_187 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_25_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_233 ();
 sky130_fd_sc_hs__fill_4 FILLER_25_241 ();
 sky130_fd_sc_hs__fill_1 FILLER_25_245 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_257 ();
 sky130_fd_sc_hs__fill_4 FILLER_25_265 ();
 sky130_fd_sc_hs__fill_1 FILLER_25_269 ();
 sky130_fd_sc_hs__fill_2 FILLER_25_288 ();
 sky130_fd_sc_hs__fill_4 FILLER_25_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_298 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_306 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_314 ();
 sky130_fd_sc_hs__fill_2 FILLER_25_322 ();
 sky130_fd_sc_hs__fill_1 FILLER_25_324 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_332 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_340 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_357 ();
 sky130_fd_sc_hs__fill_1 FILLER_25_365 ();
 sky130_fd_sc_hs__fill_4 FILLER_25_371 ();
 sky130_fd_sc_hs__fill_2 FILLER_25_375 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_398 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_25_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_25_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_25_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_25_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_26_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_26_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_26_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_88 ();
 sky130_fd_sc_hs__fill_4 FILLER_26_102 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_109 ();
 sky130_fd_sc_hs__fill_4 FILLER_26_117 ();
 sky130_fd_sc_hs__fill_2 FILLER_26_121 ();
 sky130_fd_sc_hs__fill_1 FILLER_26_126 ();
 sky130_fd_sc_hs__fill_4 FILLER_26_138 ();
 sky130_fd_sc_hs__fill_2 FILLER_26_142 ();
 sky130_fd_sc_hs__fill_1 FILLER_26_144 ();
 sky130_fd_sc_hs__fill_4 FILLER_26_146 ();
 sky130_fd_sc_hs__fill_4 FILLER_26_156 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_26_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_26_260 ();
 sky130_fd_sc_hs__fill_1 FILLER_26_262 ();
 sky130_fd_sc_hs__fill_2 FILLER_26_282 ();
 sky130_fd_sc_hs__fill_2 FILLER_26_291 ();
 sky130_fd_sc_hs__fill_1 FILLER_26_293 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_307 ();
 sky130_fd_sc_hs__fill_4 FILLER_26_315 ();
 sky130_fd_sc_hs__fill_4 FILLER_26_356 ();
 sky130_fd_sc_hs__fill_2 FILLER_26_360 ();
 sky130_fd_sc_hs__fill_4 FILLER_26_369 ();
 sky130_fd_sc_hs__fill_1 FILLER_26_376 ();
 sky130_fd_sc_hs__fill_4 FILLER_26_378 ();
 sky130_fd_sc_hs__fill_1 FILLER_26_382 ();
 sky130_fd_sc_hs__fill_2 FILLER_26_386 ();
 sky130_fd_sc_hs__fill_1 FILLER_26_388 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_413 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_421 ();
 sky130_fd_sc_hs__fill_4 FILLER_26_429 ();
 sky130_fd_sc_hs__fill_2 FILLER_26_433 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_26_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_26_526 ();
 sky130_fd_sc_hs__fill_4 FILLER_26_534 ();
 sky130_fd_sc_hs__fill_2 FILLER_26_538 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_0 ();
 sky130_fd_sc_hs__fill_4 FILLER_27_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_20 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_36 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_44 ();
 sky130_fd_sc_hs__fill_4 FILLER_27_52 ();
 sky130_fd_sc_hs__fill_2 FILLER_27_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_67 ();
 sky130_fd_sc_hs__fill_4 FILLER_27_75 ();
 sky130_fd_sc_hs__fill_1 FILLER_27_79 ();
 sky130_fd_sc_hs__fill_1 FILLER_27_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_105 ();
 sky130_fd_sc_hs__fill_2 FILLER_27_117 ();
 sky130_fd_sc_hs__fill_2 FILLER_27_130 ();
 sky130_fd_sc_hs__fill_1 FILLER_27_132 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_138 ();
 sky130_fd_sc_hs__fill_2 FILLER_27_146 ();
 sky130_fd_sc_hs__fill_2 FILLER_27_158 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_163 ();
 sky130_fd_sc_hs__fill_2 FILLER_27_171 ();
 sky130_fd_sc_hs__fill_1 FILLER_27_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_193 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_201 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_209 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_217 ();
 sky130_fd_sc_hs__fill_4 FILLER_27_225 ();
 sky130_fd_sc_hs__fill_2 FILLER_27_229 ();
 sky130_fd_sc_hs__fill_1 FILLER_27_231 ();
 sky130_fd_sc_hs__fill_4 FILLER_27_233 ();
 sky130_fd_sc_hs__fill_1 FILLER_27_237 ();
 sky130_fd_sc_hs__fill_2 FILLER_27_243 ();
 sky130_fd_sc_hs__fill_1 FILLER_27_245 ();
 sky130_fd_sc_hs__fill_4 FILLER_27_267 ();
 sky130_fd_sc_hs__fill_2 FILLER_27_271 ();
 sky130_fd_sc_hs__fill_4 FILLER_27_280 ();
 sky130_fd_sc_hs__fill_2 FILLER_27_284 ();
 sky130_fd_sc_hs__fill_1 FILLER_27_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_310 ();
 sky130_fd_sc_hs__fill_2 FILLER_27_318 ();
 sky130_fd_sc_hs__fill_1 FILLER_27_320 ();
 sky130_fd_sc_hs__fill_1 FILLER_27_324 ();
 sky130_fd_sc_hs__fill_4 FILLER_27_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_335 ();
 sky130_fd_sc_hs__fill_4 FILLER_27_343 ();
 sky130_fd_sc_hs__fill_1 FILLER_27_347 ();
 sky130_fd_sc_hs__fill_4 FILLER_27_349 ();
 sky130_fd_sc_hs__fill_2 FILLER_27_353 ();
 sky130_fd_sc_hs__fill_4 FILLER_27_358 ();
 sky130_fd_sc_hs__fill_2 FILLER_27_362 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_367 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_375 ();
 sky130_fd_sc_hs__fill_4 FILLER_27_383 ();
 sky130_fd_sc_hs__fill_2 FILLER_27_387 ();
 sky130_fd_sc_hs__fill_4 FILLER_27_399 ();
 sky130_fd_sc_hs__fill_2 FILLER_27_403 ();
 sky130_fd_sc_hs__fill_1 FILLER_27_405 ();
 sky130_fd_sc_hs__fill_1 FILLER_27_407 ();
 sky130_fd_sc_hs__fill_4 FILLER_27_411 ();
 sky130_fd_sc_hs__fill_1 FILLER_27_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_419 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_427 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_435 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_443 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_451 ();
 sky130_fd_sc_hs__fill_4 FILLER_27_459 ();
 sky130_fd_sc_hs__fill_1 FILLER_27_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_27_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_27_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_27_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_0 ();
 sky130_fd_sc_hs__fill_1 FILLER_28_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_17 ();
 sky130_fd_sc_hs__fill_4 FILLER_28_25 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_28_86 ();
 sky130_fd_sc_hs__fill_1 FILLER_28_88 ();
 sky130_fd_sc_hs__fill_4 FILLER_28_95 ();
 sky130_fd_sc_hs__fill_2 FILLER_28_99 ();
 sky130_fd_sc_hs__fill_1 FILLER_28_101 ();
 sky130_fd_sc_hs__fill_4 FILLER_28_120 ();
 sky130_fd_sc_hs__fill_4 FILLER_28_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_168 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_176 ();
 sky130_fd_sc_hs__fill_1 FILLER_28_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_212 ();
 sky130_fd_sc_hs__fill_1 FILLER_28_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_239 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_247 ();
 sky130_fd_sc_hs__fill_4 FILLER_28_255 ();
 sky130_fd_sc_hs__fill_2 FILLER_28_259 ();
 sky130_fd_sc_hs__fill_2 FILLER_28_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_271 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_279 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_287 ();
 sky130_fd_sc_hs__fill_1 FILLER_28_295 ();
 sky130_fd_sc_hs__fill_4 FILLER_28_314 ();
 sky130_fd_sc_hs__fill_1 FILLER_28_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_338 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_346 ();
 sky130_fd_sc_hs__fill_4 FILLER_28_354 ();
 sky130_fd_sc_hs__fill_1 FILLER_28_358 ();
 sky130_fd_sc_hs__fill_2 FILLER_28_378 ();
 sky130_fd_sc_hs__fill_1 FILLER_28_380 ();
 sky130_fd_sc_hs__fill_4 FILLER_28_384 ();
 sky130_fd_sc_hs__fill_1 FILLER_28_388 ();
 sky130_fd_sc_hs__fill_4 FILLER_28_394 ();
 sky130_fd_sc_hs__fill_2 FILLER_28_398 ();
 sky130_fd_sc_hs__fill_1 FILLER_28_403 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_422 ();
 sky130_fd_sc_hs__fill_4 FILLER_28_430 ();
 sky130_fd_sc_hs__fill_1 FILLER_28_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_28_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_28_526 ();
 sky130_fd_sc_hs__fill_4 FILLER_28_534 ();
 sky130_fd_sc_hs__fill_2 FILLER_28_538 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_29_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_29_115 ();
 sky130_fd_sc_hs__fill_2 FILLER_29_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_122 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_130 ();
 sky130_fd_sc_hs__fill_2 FILLER_29_138 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_153 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_161 ();
 sky130_fd_sc_hs__fill_4 FILLER_29_169 ();
 sky130_fd_sc_hs__fill_1 FILLER_29_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_199 ();
 sky130_fd_sc_hs__fill_2 FILLER_29_207 ();
 sky130_fd_sc_hs__fill_4 FILLER_29_227 ();
 sky130_fd_sc_hs__fill_1 FILLER_29_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_241 ();
 sky130_fd_sc_hs__fill_2 FILLER_29_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_258 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_266 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_274 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_282 ();
 sky130_fd_sc_hs__fill_4 FILLER_29_291 ();
 sky130_fd_sc_hs__fill_1 FILLER_29_295 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_302 ();
 sky130_fd_sc_hs__fill_1 FILLER_29_310 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_330 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_338 ();
 sky130_fd_sc_hs__fill_2 FILLER_29_346 ();
 sky130_fd_sc_hs__fill_1 FILLER_29_349 ();
 sky130_fd_sc_hs__fill_4 FILLER_29_361 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_368 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_384 ();
 sky130_fd_sc_hs__fill_4 FILLER_29_392 ();
 sky130_fd_sc_hs__fill_1 FILLER_29_396 ();
 sky130_fd_sc_hs__fill_2 FILLER_29_400 ();
 sky130_fd_sc_hs__fill_1 FILLER_29_402 ();
 sky130_fd_sc_hs__fill_2 FILLER_29_407 ();
 sky130_fd_sc_hs__fill_1 FILLER_29_409 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_413 ();
 sky130_fd_sc_hs__fill_4 FILLER_29_421 ();
 sky130_fd_sc_hs__fill_1 FILLER_29_425 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_429 ();
 sky130_fd_sc_hs__fill_4 FILLER_29_437 ();
 sky130_fd_sc_hs__fill_1 FILLER_29_441 ();
 sky130_fd_sc_hs__fill_2 FILLER_29_445 ();
 sky130_fd_sc_hs__fill_1 FILLER_29_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_451 ();
 sky130_fd_sc_hs__fill_4 FILLER_29_459 ();
 sky130_fd_sc_hs__fill_1 FILLER_29_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_29_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_29_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_29_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_30_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_30_28 ();
 sky130_fd_sc_hs__fill_4 FILLER_30_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_42 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_50 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_58 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_66 ();
 sky130_fd_sc_hs__fill_4 FILLER_30_74 ();
 sky130_fd_sc_hs__fill_1 FILLER_30_78 ();
 sky130_fd_sc_hs__fill_4 FILLER_30_82 ();
 sky130_fd_sc_hs__fill_1 FILLER_30_86 ();
 sky130_fd_sc_hs__fill_2 FILLER_30_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_96 ();
 sky130_fd_sc_hs__fill_4 FILLER_30_104 ();
 sky130_fd_sc_hs__fill_2 FILLER_30_108 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_123 ();
 sky130_fd_sc_hs__fill_2 FILLER_30_131 ();
 sky130_fd_sc_hs__fill_1 FILLER_30_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_30_202 ();
 sky130_fd_sc_hs__fill_4 FILLER_30_204 ();
 sky130_fd_sc_hs__fill_2 FILLER_30_208 ();
 sky130_fd_sc_hs__fill_1 FILLER_30_210 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_249 ();
 sky130_fd_sc_hs__fill_4 FILLER_30_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_262 ();
 sky130_fd_sc_hs__fill_4 FILLER_30_270 ();
 sky130_fd_sc_hs__fill_2 FILLER_30_274 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_297 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_305 ();
 sky130_fd_sc_hs__fill_4 FILLER_30_313 ();
 sky130_fd_sc_hs__fill_2 FILLER_30_317 ();
 sky130_fd_sc_hs__fill_2 FILLER_30_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_328 ();
 sky130_fd_sc_hs__fill_2 FILLER_30_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_30_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_378 ();
 sky130_fd_sc_hs__fill_4 FILLER_30_386 ();
 sky130_fd_sc_hs__fill_1 FILLER_30_390 ();
 sky130_fd_sc_hs__fill_4 FILLER_30_409 ();
 sky130_fd_sc_hs__fill_1 FILLER_30_413 ();
 sky130_fd_sc_hs__fill_2 FILLER_30_417 ();
 sky130_fd_sc_hs__fill_1 FILLER_30_419 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_425 ();
 sky130_fd_sc_hs__fill_2 FILLER_30_433 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_454 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_462 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_470 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_478 ();
 sky130_fd_sc_hs__fill_4 FILLER_30_486 ();
 sky130_fd_sc_hs__fill_2 FILLER_30_490 ();
 sky130_fd_sc_hs__fill_1 FILLER_30_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_30_526 ();
 sky130_fd_sc_hs__fill_4 FILLER_30_534 ();
 sky130_fd_sc_hs__fill_2 FILLER_30_538 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_31_56 ();
 sky130_fd_sc_hs__fill_4 FILLER_31_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_99 ();
 sky130_fd_sc_hs__fill_2 FILLER_31_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_31_109 ();
 sky130_fd_sc_hs__fill_1 FILLER_31_115 ();
 sky130_fd_sc_hs__fill_1 FILLER_31_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_126 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_134 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_142 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_150 ();
 sky130_fd_sc_hs__fill_1 FILLER_31_158 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_162 ();
 sky130_fd_sc_hs__fill_4 FILLER_31_170 ();
 sky130_fd_sc_hs__fill_2 FILLER_31_175 ();
 sky130_fd_sc_hs__fill_1 FILLER_31_177 ();
 sky130_fd_sc_hs__fill_1 FILLER_31_224 ();
 sky130_fd_sc_hs__fill_2 FILLER_31_230 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_241 ();
 sky130_fd_sc_hs__fill_2 FILLER_31_249 ();
 sky130_fd_sc_hs__fill_1 FILLER_31_251 ();
 sky130_fd_sc_hs__fill_4 FILLER_31_255 ();
 sky130_fd_sc_hs__fill_1 FILLER_31_259 ();
 sky130_fd_sc_hs__fill_1 FILLER_31_265 ();
 sky130_fd_sc_hs__fill_4 FILLER_31_320 ();
 sky130_fd_sc_hs__fill_2 FILLER_31_324 ();
 sky130_fd_sc_hs__fill_1 FILLER_31_326 ();
 sky130_fd_sc_hs__fill_4 FILLER_31_332 ();
 sky130_fd_sc_hs__fill_1 FILLER_31_336 ();
 sky130_fd_sc_hs__fill_1 FILLER_31_340 ();
 sky130_fd_sc_hs__fill_4 FILLER_31_367 ();
 sky130_fd_sc_hs__fill_4 FILLER_31_389 ();
 sky130_fd_sc_hs__fill_2 FILLER_31_393 ();
 sky130_fd_sc_hs__fill_1 FILLER_31_395 ();
 sky130_fd_sc_hs__fill_4 FILLER_31_399 ();
 sky130_fd_sc_hs__fill_2 FILLER_31_403 ();
 sky130_fd_sc_hs__fill_1 FILLER_31_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_415 ();
 sky130_fd_sc_hs__fill_4 FILLER_31_423 ();
 sky130_fd_sc_hs__fill_2 FILLER_31_427 ();
 sky130_fd_sc_hs__fill_1 FILLER_31_450 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_454 ();
 sky130_fd_sc_hs__fill_2 FILLER_31_462 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_31_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_31_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_31_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_32_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_32_28 ();
 sky130_fd_sc_hs__fill_1 FILLER_32_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_39 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_47 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_55 ();
 sky130_fd_sc_hs__fill_2 FILLER_32_63 ();
 sky130_fd_sc_hs__fill_1 FILLER_32_65 ();
 sky130_fd_sc_hs__fill_2 FILLER_32_85 ();
 sky130_fd_sc_hs__fill_4 FILLER_32_88 ();
 sky130_fd_sc_hs__fill_2 FILLER_32_95 ();
 sky130_fd_sc_hs__fill_1 FILLER_32_97 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_101 ();
 sky130_fd_sc_hs__fill_2 FILLER_32_109 ();
 sky130_fd_sc_hs__fill_1 FILLER_32_111 ();
 sky130_fd_sc_hs__fill_4 FILLER_32_130 ();
 sky130_fd_sc_hs__fill_1 FILLER_32_134 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_154 ();
 sky130_fd_sc_hs__fill_4 FILLER_32_162 ();
 sky130_fd_sc_hs__fill_4 FILLER_32_169 ();
 sky130_fd_sc_hs__fill_1 FILLER_32_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_192 ();
 sky130_fd_sc_hs__fill_2 FILLER_32_200 ();
 sky130_fd_sc_hs__fill_1 FILLER_32_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_222 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_230 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_238 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_246 ();
 sky130_fd_sc_hs__fill_4 FILLER_32_254 ();
 sky130_fd_sc_hs__fill_2 FILLER_32_258 ();
 sky130_fd_sc_hs__fill_1 FILLER_32_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_294 ();
 sky130_fd_sc_hs__fill_2 FILLER_32_302 ();
 sky130_fd_sc_hs__fill_1 FILLER_32_304 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_308 ();
 sky130_fd_sc_hs__fill_2 FILLER_32_316 ();
 sky130_fd_sc_hs__fill_1 FILLER_32_318 ();
 sky130_fd_sc_hs__fill_4 FILLER_32_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_342 ();
 sky130_fd_sc_hs__fill_2 FILLER_32_350 ();
 sky130_fd_sc_hs__fill_4 FILLER_32_355 ();
 sky130_fd_sc_hs__fill_1 FILLER_32_359 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_363 ();
 sky130_fd_sc_hs__fill_2 FILLER_32_371 ();
 sky130_fd_sc_hs__fill_1 FILLER_32_376 ();
 sky130_fd_sc_hs__fill_4 FILLER_32_378 ();
 sky130_fd_sc_hs__fill_2 FILLER_32_382 ();
 sky130_fd_sc_hs__fill_1 FILLER_32_384 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_388 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_396 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_404 ();
 sky130_fd_sc_hs__fill_4 FILLER_32_412 ();
 sky130_fd_sc_hs__fill_1 FILLER_32_416 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_420 ();
 sky130_fd_sc_hs__fill_4 FILLER_32_428 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_32_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_32_526 ();
 sky130_fd_sc_hs__fill_4 FILLER_32_534 ();
 sky130_fd_sc_hs__fill_2 FILLER_32_538 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_8 ();
 sky130_fd_sc_hs__fill_4 FILLER_33_16 ();
 sky130_fd_sc_hs__fill_2 FILLER_33_20 ();
 sky130_fd_sc_hs__fill_1 FILLER_33_22 ();
 sky130_fd_sc_hs__fill_2 FILLER_33_31 ();
 sky130_fd_sc_hs__fill_1 FILLER_33_33 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_42 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_50 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_59 ();
 sky130_fd_sc_hs__fill_4 FILLER_33_67 ();
 sky130_fd_sc_hs__fill_2 FILLER_33_74 ();
 sky130_fd_sc_hs__fill_2 FILLER_33_79 ();
 sky130_fd_sc_hs__fill_1 FILLER_33_81 ();
 sky130_fd_sc_hs__fill_2 FILLER_33_85 ();
 sky130_fd_sc_hs__fill_1 FILLER_33_87 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_33_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_125 ();
 sky130_fd_sc_hs__fill_2 FILLER_33_133 ();
 sky130_fd_sc_hs__fill_1 FILLER_33_135 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_147 ();
 sky130_fd_sc_hs__fill_1 FILLER_33_155 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_175 ();
 sky130_fd_sc_hs__fill_4 FILLER_33_183 ();
 sky130_fd_sc_hs__fill_1 FILLER_33_201 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_205 ();
 sky130_fd_sc_hs__fill_4 FILLER_33_213 ();
 sky130_fd_sc_hs__fill_2 FILLER_33_217 ();
 sky130_fd_sc_hs__fill_1 FILLER_33_219 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_33_231 ();
 sky130_fd_sc_hs__fill_4 FILLER_33_233 ();
 sky130_fd_sc_hs__fill_2 FILLER_33_237 ();
 sky130_fd_sc_hs__fill_1 FILLER_33_239 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_259 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_267 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_275 ();
 sky130_fd_sc_hs__fill_4 FILLER_33_283 ();
 sky130_fd_sc_hs__fill_2 FILLER_33_287 ();
 sky130_fd_sc_hs__fill_1 FILLER_33_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_307 ();
 sky130_fd_sc_hs__fill_4 FILLER_33_315 ();
 sky130_fd_sc_hs__fill_2 FILLER_33_319 ();
 sky130_fd_sc_hs__fill_1 FILLER_33_321 ();
 sky130_fd_sc_hs__fill_1 FILLER_33_329 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_333 ();
 sky130_fd_sc_hs__fill_4 FILLER_33_341 ();
 sky130_fd_sc_hs__fill_2 FILLER_33_345 ();
 sky130_fd_sc_hs__fill_1 FILLER_33_347 ();
 sky130_fd_sc_hs__fill_4 FILLER_33_372 ();
 sky130_fd_sc_hs__fill_1 FILLER_33_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_380 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_388 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_396 ();
 sky130_fd_sc_hs__fill_2 FILLER_33_404 ();
 sky130_fd_sc_hs__fill_4 FILLER_33_407 ();
 sky130_fd_sc_hs__fill_1 FILLER_33_411 ();
 sky130_fd_sc_hs__fill_2 FILLER_33_425 ();
 sky130_fd_sc_hs__fill_1 FILLER_33_427 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_33_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_33_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_33_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_33_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_34_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_34_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_54 ();
 sky130_fd_sc_hs__fill_4 FILLER_34_62 ();
 sky130_fd_sc_hs__fill_2 FILLER_34_66 ();
 sky130_fd_sc_hs__fill_1 FILLER_34_68 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_72 ();
 sky130_fd_sc_hs__fill_4 FILLER_34_80 ();
 sky130_fd_sc_hs__fill_2 FILLER_34_84 ();
 sky130_fd_sc_hs__fill_1 FILLER_34_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_104 ();
 sky130_fd_sc_hs__fill_4 FILLER_34_112 ();
 sky130_fd_sc_hs__fill_2 FILLER_34_116 ();
 sky130_fd_sc_hs__fill_4 FILLER_34_121 ();
 sky130_fd_sc_hs__fill_2 FILLER_34_125 ();
 sky130_fd_sc_hs__fill_1 FILLER_34_127 ();
 sky130_fd_sc_hs__fill_4 FILLER_34_131 ();
 sky130_fd_sc_hs__fill_4 FILLER_34_138 ();
 sky130_fd_sc_hs__fill_2 FILLER_34_142 ();
 sky130_fd_sc_hs__fill_1 FILLER_34_144 ();
 sky130_fd_sc_hs__fill_4 FILLER_34_146 ();
 sky130_fd_sc_hs__fill_1 FILLER_34_150 ();
 sky130_fd_sc_hs__fill_2 FILLER_34_172 ();
 sky130_fd_sc_hs__fill_1 FILLER_34_174 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_34_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_34_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_302 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_310 ();
 sky130_fd_sc_hs__fill_1 FILLER_34_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_344 ();
 sky130_fd_sc_hs__fill_4 FILLER_34_352 ();
 sky130_fd_sc_hs__fill_2 FILLER_34_356 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_386 ();
 sky130_fd_sc_hs__fill_2 FILLER_34_394 ();
 sky130_fd_sc_hs__fill_2 FILLER_34_414 ();
 sky130_fd_sc_hs__fill_1 FILLER_34_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_436 ();
 sky130_fd_sc_hs__fill_4 FILLER_34_447 ();
 sky130_fd_sc_hs__fill_1 FILLER_34_451 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_457 ();
 sky130_fd_sc_hs__fill_4 FILLER_34_465 ();
 sky130_fd_sc_hs__fill_1 FILLER_34_469 ();
 sky130_fd_sc_hs__fill_2 FILLER_34_473 ();
 sky130_fd_sc_hs__fill_1 FILLER_34_475 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_479 ();
 sky130_fd_sc_hs__fill_4 FILLER_34_487 ();
 sky130_fd_sc_hs__fill_2 FILLER_34_491 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_502 ();
 sky130_fd_sc_hs__fill_1 FILLER_34_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_519 ();
 sky130_fd_sc_hs__fill_8 FILLER_34_527 ();
 sky130_fd_sc_hs__fill_4 FILLER_34_535 ();
 sky130_fd_sc_hs__fill_1 FILLER_34_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_35_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_91 ();
 sky130_fd_sc_hs__fill_2 FILLER_35_99 ();
 sky130_fd_sc_hs__fill_1 FILLER_35_101 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_108 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_117 ();
 sky130_fd_sc_hs__fill_4 FILLER_35_125 ();
 sky130_fd_sc_hs__fill_2 FILLER_35_129 ();
 sky130_fd_sc_hs__fill_4 FILLER_35_168 ();
 sky130_fd_sc_hs__fill_2 FILLER_35_172 ();
 sky130_fd_sc_hs__fill_4 FILLER_35_175 ();
 sky130_fd_sc_hs__fill_1 FILLER_35_179 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_185 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_193 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_201 ();
 sky130_fd_sc_hs__fill_4 FILLER_35_209 ();
 sky130_fd_sc_hs__fill_1 FILLER_35_213 ();
 sky130_fd_sc_hs__fill_2 FILLER_35_233 ();
 sky130_fd_sc_hs__fill_1 FILLER_35_235 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_254 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_278 ();
 sky130_fd_sc_hs__fill_4 FILLER_35_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_35_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_349 ();
 sky130_fd_sc_hs__fill_2 FILLER_35_357 ();
 sky130_fd_sc_hs__fill_4 FILLER_35_362 ();
 sky130_fd_sc_hs__fill_1 FILLER_35_366 ();
 sky130_fd_sc_hs__fill_1 FILLER_35_370 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_35_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_431 ();
 sky130_fd_sc_hs__fill_4 FILLER_35_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_483 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_491 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_499 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_507 ();
 sky130_fd_sc_hs__fill_4 FILLER_35_515 ();
 sky130_fd_sc_hs__fill_2 FILLER_35_519 ();
 sky130_fd_sc_hs__fill_1 FILLER_35_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_35_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_35_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_8 ();
 sky130_fd_sc_hs__fill_4 FILLER_36_16 ();
 sky130_fd_sc_hs__fill_1 FILLER_36_20 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_73 ();
 sky130_fd_sc_hs__fill_2 FILLER_36_84 ();
 sky130_fd_sc_hs__fill_1 FILLER_36_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_96 ();
 sky130_fd_sc_hs__fill_2 FILLER_36_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_133 ();
 sky130_fd_sc_hs__fill_4 FILLER_36_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_36_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_212 ();
 sky130_fd_sc_hs__fill_4 FILLER_36_239 ();
 sky130_fd_sc_hs__fill_1 FILLER_36_243 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_247 ();
 sky130_fd_sc_hs__fill_4 FILLER_36_255 ();
 sky130_fd_sc_hs__fill_2 FILLER_36_259 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_262 ();
 sky130_fd_sc_hs__fill_4 FILLER_36_270 ();
 sky130_fd_sc_hs__fill_2 FILLER_36_274 ();
 sky130_fd_sc_hs__fill_1 FILLER_36_276 ();
 sky130_fd_sc_hs__fill_1 FILLER_36_301 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_305 ();
 sky130_fd_sc_hs__fill_2 FILLER_36_316 ();
 sky130_fd_sc_hs__fill_1 FILLER_36_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_36_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_386 ();
 sky130_fd_sc_hs__fill_1 FILLER_36_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_398 ();
 sky130_fd_sc_hs__fill_4 FILLER_36_406 ();
 sky130_fd_sc_hs__fill_1 FILLER_36_410 ();
 sky130_fd_sc_hs__fill_4 FILLER_36_414 ();
 sky130_fd_sc_hs__fill_2 FILLER_36_418 ();
 sky130_fd_sc_hs__fill_1 FILLER_36_420 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_424 ();
 sky130_fd_sc_hs__fill_2 FILLER_36_432 ();
 sky130_fd_sc_hs__fill_1 FILLER_36_434 ();
 sky130_fd_sc_hs__fill_4 FILLER_36_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_453 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_467 ();
 sky130_fd_sc_hs__fill_4 FILLER_36_475 ();
 sky130_fd_sc_hs__fill_2 FILLER_36_479 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_36_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_502 ();
 sky130_fd_sc_hs__fill_4 FILLER_36_510 ();
 sky130_fd_sc_hs__fill_2 FILLER_36_514 ();
 sky130_fd_sc_hs__fill_1 FILLER_36_516 ();
 sky130_fd_sc_hs__fill_8 FILLER_36_525 ();
 sky130_fd_sc_hs__fill_4 FILLER_36_533 ();
 sky130_fd_sc_hs__fill_2 FILLER_36_537 ();
 sky130_fd_sc_hs__fill_1 FILLER_36_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_0 ();
 sky130_fd_sc_hs__fill_2 FILLER_37_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_18 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_26 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_34 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_42 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_50 ();
 sky130_fd_sc_hs__fill_4 FILLER_37_59 ();
 sky130_fd_sc_hs__fill_2 FILLER_37_63 ();
 sky130_fd_sc_hs__fill_1 FILLER_37_65 ();
 sky130_fd_sc_hs__fill_4 FILLER_37_75 ();
 sky130_fd_sc_hs__fill_1 FILLER_37_97 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_37_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_215 ();
 sky130_fd_sc_hs__fill_2 FILLER_37_223 ();
 sky130_fd_sc_hs__fill_4 FILLER_37_228 ();
 sky130_fd_sc_hs__fill_2 FILLER_37_233 ();
 sky130_fd_sc_hs__fill_2 FILLER_37_259 ();
 sky130_fd_sc_hs__fill_1 FILLER_37_261 ();
 sky130_fd_sc_hs__fill_1 FILLER_37_286 ();
 sky130_fd_sc_hs__fill_4 FILLER_37_337 ();
 sky130_fd_sc_hs__fill_1 FILLER_37_341 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_365 ();
 sky130_fd_sc_hs__fill_2 FILLER_37_373 ();
 sky130_fd_sc_hs__fill_1 FILLER_37_375 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_379 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_387 ();
 sky130_fd_sc_hs__fill_4 FILLER_37_395 ();
 sky130_fd_sc_hs__fill_1 FILLER_37_405 ();
 sky130_fd_sc_hs__fill_4 FILLER_37_407 ();
 sky130_fd_sc_hs__fill_2 FILLER_37_411 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_442 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_450 ();
 sky130_fd_sc_hs__fill_4 FILLER_37_458 ();
 sky130_fd_sc_hs__fill_2 FILLER_37_462 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_497 ();
 sky130_fd_sc_hs__fill_1 FILLER_37_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_514 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_37_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_37_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_38_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_38_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_46 ();
 sky130_fd_sc_hs__fill_1 FILLER_38_54 ();
 sky130_fd_sc_hs__fill_2 FILLER_38_67 ();
 sky130_fd_sc_hs__fill_1 FILLER_38_69 ();
 sky130_fd_sc_hs__fill_4 FILLER_38_73 ();
 sky130_fd_sc_hs__fill_4 FILLER_38_80 ();
 sky130_fd_sc_hs__fill_2 FILLER_38_84 ();
 sky130_fd_sc_hs__fill_1 FILLER_38_86 ();
 sky130_fd_sc_hs__fill_1 FILLER_38_91 ();
 sky130_fd_sc_hs__fill_4 FILLER_38_95 ();
 sky130_fd_sc_hs__fill_1 FILLER_38_102 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_162 ();
 sky130_fd_sc_hs__fill_2 FILLER_38_170 ();
 sky130_fd_sc_hs__fill_4 FILLER_38_179 ();
 sky130_fd_sc_hs__fill_1 FILLER_38_183 ();
 sky130_fd_sc_hs__fill_1 FILLER_38_187 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_38_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_204 ();
 sky130_fd_sc_hs__fill_2 FILLER_38_212 ();
 sky130_fd_sc_hs__fill_2 FILLER_38_217 ();
 sky130_fd_sc_hs__fill_1 FILLER_38_219 ();
 sky130_fd_sc_hs__fill_4 FILLER_38_223 ();
 sky130_fd_sc_hs__fill_2 FILLER_38_227 ();
 sky130_fd_sc_hs__fill_4 FILLER_38_232 ();
 sky130_fd_sc_hs__fill_4 FILLER_38_257 ();
 sky130_fd_sc_hs__fill_1 FILLER_38_262 ();
 sky130_fd_sc_hs__fill_1 FILLER_38_269 ();
 sky130_fd_sc_hs__fill_2 FILLER_38_291 ();
 sky130_fd_sc_hs__fill_4 FILLER_38_296 ();
 sky130_fd_sc_hs__fill_4 FILLER_38_323 ();
 sky130_fd_sc_hs__fill_1 FILLER_38_330 ();
 sky130_fd_sc_hs__fill_1 FILLER_38_350 ();
 sky130_fd_sc_hs__fill_2 FILLER_38_354 ();
 sky130_fd_sc_hs__fill_2 FILLER_38_374 ();
 sky130_fd_sc_hs__fill_1 FILLER_38_376 ();
 sky130_fd_sc_hs__fill_2 FILLER_38_378 ();
 sky130_fd_sc_hs__fill_1 FILLER_38_380 ();
 sky130_fd_sc_hs__fill_1 FILLER_38_384 ();
 sky130_fd_sc_hs__fill_1 FILLER_38_404 ();
 sky130_fd_sc_hs__fill_1 FILLER_38_423 ();
 sky130_fd_sc_hs__fill_2 FILLER_38_427 ();
 sky130_fd_sc_hs__fill_2 FILLER_38_432 ();
 sky130_fd_sc_hs__fill_1 FILLER_38_434 ();
 sky130_fd_sc_hs__fill_2 FILLER_38_439 ();
 sky130_fd_sc_hs__fill_1 FILLER_38_441 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_445 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_453 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_461 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_469 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_477 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_485 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_494 ();
 sky130_fd_sc_hs__fill_1 FILLER_38_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_511 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_519 ();
 sky130_fd_sc_hs__fill_8 FILLER_38_527 ();
 sky130_fd_sc_hs__fill_4 FILLER_38_535 ();
 sky130_fd_sc_hs__fill_1 FILLER_38_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_8 ();
 sky130_fd_sc_hs__fill_2 FILLER_39_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_34 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_42 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_50 ();
 sky130_fd_sc_hs__fill_4 FILLER_39_59 ();
 sky130_fd_sc_hs__fill_2 FILLER_39_63 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_86 ();
 sky130_fd_sc_hs__fill_4 FILLER_39_94 ();
 sky130_fd_sc_hs__fill_2 FILLER_39_98 ();
 sky130_fd_sc_hs__fill_1 FILLER_39_100 ();
 sky130_fd_sc_hs__fill_2 FILLER_39_104 ();
 sky130_fd_sc_hs__fill_1 FILLER_39_106 ();
 sky130_fd_sc_hs__fill_2 FILLER_39_110 ();
 sky130_fd_sc_hs__fill_1 FILLER_39_115 ();
 sky130_fd_sc_hs__fill_1 FILLER_39_120 ();
 sky130_fd_sc_hs__fill_2 FILLER_39_124 ();
 sky130_fd_sc_hs__fill_1 FILLER_39_126 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_130 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_138 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_162 ();
 sky130_fd_sc_hs__fill_4 FILLER_39_170 ();
 sky130_fd_sc_hs__fill_4 FILLER_39_175 ();
 sky130_fd_sc_hs__fill_1 FILLER_39_179 ();
 sky130_fd_sc_hs__fill_2 FILLER_39_198 ();
 sky130_fd_sc_hs__fill_2 FILLER_39_206 ();
 sky130_fd_sc_hs__fill_1 FILLER_39_208 ();
 sky130_fd_sc_hs__fill_4 FILLER_39_227 ();
 sky130_fd_sc_hs__fill_1 FILLER_39_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_252 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_268 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_276 ();
 sky130_fd_sc_hs__fill_4 FILLER_39_284 ();
 sky130_fd_sc_hs__fill_2 FILLER_39_288 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_307 ();
 sky130_fd_sc_hs__fill_1 FILLER_39_315 ();
 sky130_fd_sc_hs__fill_1 FILLER_39_340 ();
 sky130_fd_sc_hs__fill_2 FILLER_39_346 ();
 sky130_fd_sc_hs__fill_2 FILLER_39_370 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_393 ();
 sky130_fd_sc_hs__fill_4 FILLER_39_401 ();
 sky130_fd_sc_hs__fill_1 FILLER_39_405 ();
 sky130_fd_sc_hs__fill_2 FILLER_39_407 ();
 sky130_fd_sc_hs__fill_1 FILLER_39_409 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_39_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_39_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_39_521 ();
 sky130_fd_sc_hs__fill_4 FILLER_39_523 ();
 sky130_fd_sc_hs__fill_2 FILLER_39_527 ();
 sky130_fd_sc_hs__fill_2 FILLER_39_537 ();
 sky130_fd_sc_hs__fill_1 FILLER_39_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_40_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_40_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_73 ();
 sky130_fd_sc_hs__fill_4 FILLER_40_81 ();
 sky130_fd_sc_hs__fill_2 FILLER_40_85 ();
 sky130_fd_sc_hs__fill_4 FILLER_40_88 ();
 sky130_fd_sc_hs__fill_1 FILLER_40_92 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_111 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_119 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_127 ();
 sky130_fd_sc_hs__fill_2 FILLER_40_146 ();
 sky130_fd_sc_hs__fill_4 FILLER_40_166 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_191 ();
 sky130_fd_sc_hs__fill_4 FILLER_40_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_223 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_231 ();
 sky130_fd_sc_hs__fill_4 FILLER_40_239 ();
 sky130_fd_sc_hs__fill_2 FILLER_40_243 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_248 ();
 sky130_fd_sc_hs__fill_4 FILLER_40_256 ();
 sky130_fd_sc_hs__fill_1 FILLER_40_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_262 ();
 sky130_fd_sc_hs__fill_4 FILLER_40_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_277 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_285 ();
 sky130_fd_sc_hs__fill_2 FILLER_40_293 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_298 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_306 ();
 sky130_fd_sc_hs__fill_4 FILLER_40_314 ();
 sky130_fd_sc_hs__fill_1 FILLER_40_318 ();
 sky130_fd_sc_hs__fill_4 FILLER_40_329 ();
 sky130_fd_sc_hs__fill_1 FILLER_40_363 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_367 ();
 sky130_fd_sc_hs__fill_2 FILLER_40_375 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_410 ();
 sky130_fd_sc_hs__fill_4 FILLER_40_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_425 ();
 sky130_fd_sc_hs__fill_2 FILLER_40_433 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_436 ();
 sky130_fd_sc_hs__fill_4 FILLER_40_444 ();
 sky130_fd_sc_hs__fill_2 FILLER_40_448 ();
 sky130_fd_sc_hs__fill_1 FILLER_40_450 ();
 sky130_fd_sc_hs__fill_4 FILLER_40_454 ();
 sky130_fd_sc_hs__fill_2 FILLER_40_458 ();
 sky130_fd_sc_hs__fill_4 FILLER_40_466 ();
 sky130_fd_sc_hs__fill_4 FILLER_40_488 ();
 sky130_fd_sc_hs__fill_1 FILLER_40_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_40_526 ();
 sky130_fd_sc_hs__fill_4 FILLER_40_534 ();
 sky130_fd_sc_hs__fill_2 FILLER_40_538 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_41_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_67 ();
 sky130_fd_sc_hs__fill_1 FILLER_41_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_79 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_87 ();
 sky130_fd_sc_hs__fill_4 FILLER_41_95 ();
 sky130_fd_sc_hs__fill_1 FILLER_41_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_103 ();
 sky130_fd_sc_hs__fill_4 FILLER_41_111 ();
 sky130_fd_sc_hs__fill_1 FILLER_41_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_125 ();
 sky130_fd_sc_hs__fill_4 FILLER_41_133 ();
 sky130_fd_sc_hs__fill_2 FILLER_41_137 ();
 sky130_fd_sc_hs__fill_4 FILLER_41_164 ();
 sky130_fd_sc_hs__fill_2 FILLER_41_171 ();
 sky130_fd_sc_hs__fill_1 FILLER_41_173 ();
 sky130_fd_sc_hs__fill_1 FILLER_41_193 ();
 sky130_fd_sc_hs__fill_2 FILLER_41_212 ();
 sky130_fd_sc_hs__fill_1 FILLER_41_214 ();
 sky130_fd_sc_hs__fill_2 FILLER_41_218 ();
 sky130_fd_sc_hs__fill_1 FILLER_41_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_224 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_251 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_259 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_270 ();
 sky130_fd_sc_hs__fill_4 FILLER_41_278 ();
 sky130_fd_sc_hs__fill_2 FILLER_41_282 ();
 sky130_fd_sc_hs__fill_1 FILLER_41_284 ();
 sky130_fd_sc_hs__fill_2 FILLER_41_288 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_302 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_313 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_321 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_329 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_337 ();
 sky130_fd_sc_hs__fill_2 FILLER_41_345 ();
 sky130_fd_sc_hs__fill_1 FILLER_41_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_349 ();
 sky130_fd_sc_hs__fill_4 FILLER_41_357 ();
 sky130_fd_sc_hs__fill_2 FILLER_41_361 ();
 sky130_fd_sc_hs__fill_1 FILLER_41_363 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_387 ();
 sky130_fd_sc_hs__fill_4 FILLER_41_395 ();
 sky130_fd_sc_hs__fill_2 FILLER_41_399 ();
 sky130_fd_sc_hs__fill_2 FILLER_41_404 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_415 ();
 sky130_fd_sc_hs__fill_1 FILLER_41_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_427 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_435 ();
 sky130_fd_sc_hs__fill_2 FILLER_41_443 ();
 sky130_fd_sc_hs__fill_1 FILLER_41_445 ();
 sky130_fd_sc_hs__fill_4 FILLER_41_465 ();
 sky130_fd_sc_hs__fill_1 FILLER_41_469 ();
 sky130_fd_sc_hs__fill_2 FILLER_41_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_486 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_510 ();
 sky130_fd_sc_hs__fill_4 FILLER_41_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_41_523 ();
 sky130_fd_sc_hs__fill_1 FILLER_41_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_42_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_42_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_38 ();
 sky130_fd_sc_hs__fill_4 FILLER_42_46 ();
 sky130_fd_sc_hs__fill_2 FILLER_42_50 ();
 sky130_fd_sc_hs__fill_4 FILLER_42_62 ();
 sky130_fd_sc_hs__fill_2 FILLER_42_66 ();
 sky130_fd_sc_hs__fill_1 FILLER_42_68 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_120 ();
 sky130_fd_sc_hs__fill_4 FILLER_42_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_135 ();
 sky130_fd_sc_hs__fill_2 FILLER_42_143 ();
 sky130_fd_sc_hs__fill_1 FILLER_42_146 ();
 sky130_fd_sc_hs__fill_1 FILLER_42_150 ();
 sky130_fd_sc_hs__fill_2 FILLER_42_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_177 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_185 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_193 ();
 sky130_fd_sc_hs__fill_2 FILLER_42_201 ();
 sky130_fd_sc_hs__fill_4 FILLER_42_204 ();
 sky130_fd_sc_hs__fill_2 FILLER_42_208 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_213 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_221 ();
 sky130_fd_sc_hs__fill_2 FILLER_42_229 ();
 sky130_fd_sc_hs__fill_2 FILLER_42_234 ();
 sky130_fd_sc_hs__fill_1 FILLER_42_236 ();
 sky130_fd_sc_hs__fill_4 FILLER_42_240 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_247 ();
 sky130_fd_sc_hs__fill_4 FILLER_42_255 ();
 sky130_fd_sc_hs__fill_2 FILLER_42_259 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_298 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_306 ();
 sky130_fd_sc_hs__fill_4 FILLER_42_314 ();
 sky130_fd_sc_hs__fill_1 FILLER_42_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_352 ();
 sky130_fd_sc_hs__fill_1 FILLER_42_360 ();
 sky130_fd_sc_hs__fill_4 FILLER_42_370 ();
 sky130_fd_sc_hs__fill_2 FILLER_42_374 ();
 sky130_fd_sc_hs__fill_1 FILLER_42_376 ();
 sky130_fd_sc_hs__fill_1 FILLER_42_378 ();
 sky130_fd_sc_hs__fill_4 FILLER_42_386 ();
 sky130_fd_sc_hs__fill_2 FILLER_42_390 ();
 sky130_fd_sc_hs__fill_1 FILLER_42_392 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_454 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_510 ();
 sky130_fd_sc_hs__fill_4 FILLER_42_518 ();
 sky130_fd_sc_hs__fill_2 FILLER_42_522 ();
 sky130_fd_sc_hs__fill_8 FILLER_42_532 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_43_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_59 ();
 sky130_fd_sc_hs__fill_2 FILLER_43_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_72 ();
 sky130_fd_sc_hs__fill_1 FILLER_43_80 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_43_115 ();
 sky130_fd_sc_hs__fill_4 FILLER_43_117 ();
 sky130_fd_sc_hs__fill_2 FILLER_43_139 ();
 sky130_fd_sc_hs__fill_1 FILLER_43_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_145 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_153 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_161 ();
 sky130_fd_sc_hs__fill_4 FILLER_43_169 ();
 sky130_fd_sc_hs__fill_1 FILLER_43_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_43_231 ();
 sky130_fd_sc_hs__fill_2 FILLER_43_233 ();
 sky130_fd_sc_hs__fill_1 FILLER_43_235 ();
 sky130_fd_sc_hs__fill_1 FILLER_43_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_261 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_314 ();
 sky130_fd_sc_hs__fill_1 FILLER_43_322 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_326 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_334 ();
 sky130_fd_sc_hs__fill_4 FILLER_43_342 ();
 sky130_fd_sc_hs__fill_2 FILLER_43_346 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_373 ();
 sky130_fd_sc_hs__fill_4 FILLER_43_381 ();
 sky130_fd_sc_hs__fill_1 FILLER_43_385 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_395 ();
 sky130_fd_sc_hs__fill_2 FILLER_43_403 ();
 sky130_fd_sc_hs__fill_1 FILLER_43_405 ();
 sky130_fd_sc_hs__fill_2 FILLER_43_407 ();
 sky130_fd_sc_hs__fill_1 FILLER_43_409 ();
 sky130_fd_sc_hs__fill_4 FILLER_43_419 ();
 sky130_fd_sc_hs__fill_2 FILLER_43_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_449 ();
 sky130_fd_sc_hs__fill_4 FILLER_43_457 ();
 sky130_fd_sc_hs__fill_2 FILLER_43_461 ();
 sky130_fd_sc_hs__fill_1 FILLER_43_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_473 ();
 sky130_fd_sc_hs__fill_4 FILLER_43_481 ();
 sky130_fd_sc_hs__fill_2 FILLER_43_485 ();
 sky130_fd_sc_hs__fill_1 FILLER_43_487 ();
 sky130_fd_sc_hs__fill_1 FILLER_43_491 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_495 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_503 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_511 ();
 sky130_fd_sc_hs__fill_2 FILLER_43_519 ();
 sky130_fd_sc_hs__fill_1 FILLER_43_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_43_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_43_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_0 ();
 sky130_fd_sc_hs__fill_1 FILLER_44_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_17 ();
 sky130_fd_sc_hs__fill_4 FILLER_44_25 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_46 ();
 sky130_fd_sc_hs__fill_2 FILLER_44_54 ();
 sky130_fd_sc_hs__fill_1 FILLER_44_56 ();
 sky130_fd_sc_hs__fill_1 FILLER_44_78 ();
 sky130_fd_sc_hs__fill_4 FILLER_44_82 ();
 sky130_fd_sc_hs__fill_1 FILLER_44_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_88 ();
 sky130_fd_sc_hs__fill_2 FILLER_44_96 ();
 sky130_fd_sc_hs__fill_1 FILLER_44_98 ();
 sky130_fd_sc_hs__fill_4 FILLER_44_123 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_186 ();
 sky130_fd_sc_hs__fill_1 FILLER_44_194 ();
 sky130_fd_sc_hs__fill_4 FILLER_44_198 ();
 sky130_fd_sc_hs__fill_1 FILLER_44_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_223 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_231 ();
 sky130_fd_sc_hs__fill_4 FILLER_44_239 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_302 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_310 ();
 sky130_fd_sc_hs__fill_1 FILLER_44_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_328 ();
 sky130_fd_sc_hs__fill_4 FILLER_44_336 ();
 sky130_fd_sc_hs__fill_1 FILLER_44_340 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_44_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_378 ();
 sky130_fd_sc_hs__fill_4 FILLER_44_386 ();
 sky130_fd_sc_hs__fill_2 FILLER_44_390 ();
 sky130_fd_sc_hs__fill_2 FILLER_44_397 ();
 sky130_fd_sc_hs__fill_2 FILLER_44_417 ();
 sky130_fd_sc_hs__fill_1 FILLER_44_419 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_423 ();
 sky130_fd_sc_hs__fill_1 FILLER_44_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_457 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_481 ();
 sky130_fd_sc_hs__fill_4 FILLER_44_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_510 ();
 sky130_fd_sc_hs__fill_4 FILLER_44_518 ();
 sky130_fd_sc_hs__fill_2 FILLER_44_522 ();
 sky130_fd_sc_hs__fill_8 FILLER_44_532 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_45_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_62 ();
 sky130_fd_sc_hs__fill_1 FILLER_45_70 ();
 sky130_fd_sc_hs__fill_2 FILLER_45_74 ();
 sky130_fd_sc_hs__fill_1 FILLER_45_76 ();
 sky130_fd_sc_hs__fill_2 FILLER_45_113 ();
 sky130_fd_sc_hs__fill_1 FILLER_45_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_127 ();
 sky130_fd_sc_hs__fill_2 FILLER_45_135 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_155 ();
 sky130_fd_sc_hs__fill_2 FILLER_45_163 ();
 sky130_fd_sc_hs__fill_4 FILLER_45_168 ();
 sky130_fd_sc_hs__fill_2 FILLER_45_172 ();
 sky130_fd_sc_hs__fill_4 FILLER_45_175 ();
 sky130_fd_sc_hs__fill_2 FILLER_45_179 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_184 ();
 sky130_fd_sc_hs__fill_2 FILLER_45_192 ();
 sky130_fd_sc_hs__fill_1 FILLER_45_194 ();
 sky130_fd_sc_hs__fill_2 FILLER_45_216 ();
 sky130_fd_sc_hs__fill_1 FILLER_45_218 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_222 ();
 sky130_fd_sc_hs__fill_2 FILLER_45_230 ();
 sky130_fd_sc_hs__fill_4 FILLER_45_233 ();
 sky130_fd_sc_hs__fill_1 FILLER_45_237 ();
 sky130_fd_sc_hs__fill_1 FILLER_45_256 ();
 sky130_fd_sc_hs__fill_1 FILLER_45_275 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_279 ();
 sky130_fd_sc_hs__fill_2 FILLER_45_287 ();
 sky130_fd_sc_hs__fill_1 FILLER_45_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_315 ();
 sky130_fd_sc_hs__fill_4 FILLER_45_323 ();
 sky130_fd_sc_hs__fill_1 FILLER_45_327 ();
 sky130_fd_sc_hs__fill_2 FILLER_45_346 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_45_405 ();
 sky130_fd_sc_hs__fill_2 FILLER_45_407 ();
 sky130_fd_sc_hs__fill_1 FILLER_45_409 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_422 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_430 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_438 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_446 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_454 ();
 sky130_fd_sc_hs__fill_2 FILLER_45_462 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_505 ();
 sky130_fd_sc_hs__fill_1 FILLER_45_513 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_45_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_45_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_8 ();
 sky130_fd_sc_hs__fill_4 FILLER_46_16 ();
 sky130_fd_sc_hs__fill_1 FILLER_46_20 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_38 ();
 sky130_fd_sc_hs__fill_2 FILLER_46_46 ();
 sky130_fd_sc_hs__fill_1 FILLER_46_48 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_75 ();
 sky130_fd_sc_hs__fill_4 FILLER_46_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_99 ();
 sky130_fd_sc_hs__fill_2 FILLER_46_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_46_109 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_134 ();
 sky130_fd_sc_hs__fill_2 FILLER_46_142 ();
 sky130_fd_sc_hs__fill_1 FILLER_46_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_146 ();
 sky130_fd_sc_hs__fill_4 FILLER_46_154 ();
 sky130_fd_sc_hs__fill_1 FILLER_46_158 ();
 sky130_fd_sc_hs__fill_1 FILLER_46_162 ();
 sky130_fd_sc_hs__fill_4 FILLER_46_187 ();
 sky130_fd_sc_hs__fill_2 FILLER_46_191 ();
 sky130_fd_sc_hs__fill_1 FILLER_46_193 ();
 sky130_fd_sc_hs__fill_4 FILLER_46_197 ();
 sky130_fd_sc_hs__fill_2 FILLER_46_201 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_204 ();
 sky130_fd_sc_hs__fill_1 FILLER_46_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_234 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_242 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_253 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_302 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_310 ();
 sky130_fd_sc_hs__fill_1 FILLER_46_318 ();
 sky130_fd_sc_hs__fill_2 FILLER_46_374 ();
 sky130_fd_sc_hs__fill_1 FILLER_46_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_46_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_444 ();
 sky130_fd_sc_hs__fill_2 FILLER_46_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_475 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_483 ();
 sky130_fd_sc_hs__fill_2 FILLER_46_491 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_494 ();
 sky130_fd_sc_hs__fill_1 FILLER_46_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_511 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_519 ();
 sky130_fd_sc_hs__fill_8 FILLER_46_527 ();
 sky130_fd_sc_hs__fill_4 FILLER_46_535 ();
 sky130_fd_sc_hs__fill_1 FILLER_46_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_40 ();
 sky130_fd_sc_hs__fill_2 FILLER_47_48 ();
 sky130_fd_sc_hs__fill_4 FILLER_47_53 ();
 sky130_fd_sc_hs__fill_1 FILLER_47_57 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_59 ();
 sky130_fd_sc_hs__fill_4 FILLER_47_67 ();
 sky130_fd_sc_hs__fill_2 FILLER_47_71 ();
 sky130_fd_sc_hs__fill_1 FILLER_47_73 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_77 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_85 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_93 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_101 ();
 sky130_fd_sc_hs__fill_4 FILLER_47_109 ();
 sky130_fd_sc_hs__fill_2 FILLER_47_113 ();
 sky130_fd_sc_hs__fill_1 FILLER_47_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_117 ();
 sky130_fd_sc_hs__fill_4 FILLER_47_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_147 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_155 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_163 ();
 sky130_fd_sc_hs__fill_1 FILLER_47_193 ();
 sky130_fd_sc_hs__fill_2 FILLER_47_212 ();
 sky130_fd_sc_hs__fill_2 FILLER_47_217 ();
 sky130_fd_sc_hs__fill_4 FILLER_47_222 ();
 sky130_fd_sc_hs__fill_2 FILLER_47_226 ();
 sky130_fd_sc_hs__fill_1 FILLER_47_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_257 ();
 sky130_fd_sc_hs__fill_4 FILLER_47_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_272 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_280 ();
 sky130_fd_sc_hs__fill_2 FILLER_47_288 ();
 sky130_fd_sc_hs__fill_2 FILLER_47_291 ();
 sky130_fd_sc_hs__fill_1 FILLER_47_293 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_312 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_338 ();
 sky130_fd_sc_hs__fill_2 FILLER_47_346 ();
 sky130_fd_sc_hs__fill_2 FILLER_47_349 ();
 sky130_fd_sc_hs__fill_1 FILLER_47_351 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_389 ();
 sky130_fd_sc_hs__fill_4 FILLER_47_397 ();
 sky130_fd_sc_hs__fill_2 FILLER_47_404 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_473 ();
 sky130_fd_sc_hs__fill_4 FILLER_47_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_506 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_514 ();
 sky130_fd_sc_hs__fill_8 FILLER_47_523 ();
 sky130_fd_sc_hs__fill_1 FILLER_47_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_48_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_48_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_38 ();
 sky130_fd_sc_hs__fill_1 FILLER_48_46 ();
 sky130_fd_sc_hs__fill_4 FILLER_48_65 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_128 ();
 sky130_fd_sc_hs__fill_4 FILLER_48_139 ();
 sky130_fd_sc_hs__fill_2 FILLER_48_143 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_164 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_193 ();
 sky130_fd_sc_hs__fill_2 FILLER_48_201 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_204 ();
 sky130_fd_sc_hs__fill_2 FILLER_48_212 ();
 sky130_fd_sc_hs__fill_1 FILLER_48_214 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_233 ();
 sky130_fd_sc_hs__fill_2 FILLER_48_241 ();
 sky130_fd_sc_hs__fill_1 FILLER_48_262 ();
 sky130_fd_sc_hs__fill_1 FILLER_48_266 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_285 ();
 sky130_fd_sc_hs__fill_2 FILLER_48_293 ();
 sky130_fd_sc_hs__fill_4 FILLER_48_313 ();
 sky130_fd_sc_hs__fill_2 FILLER_48_317 ();
 sky130_fd_sc_hs__fill_1 FILLER_48_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_339 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_347 ();
 sky130_fd_sc_hs__fill_2 FILLER_48_355 ();
 sky130_fd_sc_hs__fill_2 FILLER_48_375 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_397 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_413 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_421 ();
 sky130_fd_sc_hs__fill_4 FILLER_48_429 ();
 sky130_fd_sc_hs__fill_2 FILLER_48_433 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_444 ();
 sky130_fd_sc_hs__fill_2 FILLER_48_452 ();
 sky130_fd_sc_hs__fill_1 FILLER_48_454 ();
 sky130_fd_sc_hs__fill_1 FILLER_48_460 ();
 sky130_fd_sc_hs__fill_2 FILLER_48_487 ();
 sky130_fd_sc_hs__fill_1 FILLER_48_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_505 ();
 sky130_fd_sc_hs__fill_2 FILLER_48_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_48_515 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_524 ();
 sky130_fd_sc_hs__fill_8 FILLER_48_532 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_40 ();
 sky130_fd_sc_hs__fill_4 FILLER_49_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_49_52 ();
 sky130_fd_sc_hs__fill_1 FILLER_49_54 ();
 sky130_fd_sc_hs__fill_4 FILLER_49_59 ();
 sky130_fd_sc_hs__fill_2 FILLER_49_63 ();
 sky130_fd_sc_hs__fill_4 FILLER_49_86 ();
 sky130_fd_sc_hs__fill_2 FILLER_49_90 ();
 sky130_fd_sc_hs__fill_1 FILLER_49_92 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_104 ();
 sky130_fd_sc_hs__fill_4 FILLER_49_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_117 ();
 sky130_fd_sc_hs__fill_4 FILLER_49_125 ();
 sky130_fd_sc_hs__fill_2 FILLER_49_129 ();
 sky130_fd_sc_hs__fill_1 FILLER_49_131 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_153 ();
 sky130_fd_sc_hs__fill_4 FILLER_49_161 ();
 sky130_fd_sc_hs__fill_2 FILLER_49_165 ();
 sky130_fd_sc_hs__fill_2 FILLER_49_172 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_175 ();
 sky130_fd_sc_hs__fill_1 FILLER_49_183 ();
 sky130_fd_sc_hs__fill_1 FILLER_49_187 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_199 ();
 sky130_fd_sc_hs__fill_4 FILLER_49_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_214 ();
 sky130_fd_sc_hs__fill_4 FILLER_49_222 ();
 sky130_fd_sc_hs__fill_2 FILLER_49_229 ();
 sky130_fd_sc_hs__fill_1 FILLER_49_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_251 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_259 ();
 sky130_fd_sc_hs__fill_2 FILLER_49_267 ();
 sky130_fd_sc_hs__fill_2 FILLER_49_287 ();
 sky130_fd_sc_hs__fill_1 FILLER_49_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_327 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_335 ();
 sky130_fd_sc_hs__fill_4 FILLER_49_343 ();
 sky130_fd_sc_hs__fill_1 FILLER_49_347 ();
 sky130_fd_sc_hs__fill_1 FILLER_49_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_353 ();
 sky130_fd_sc_hs__fill_1 FILLER_49_361 ();
 sky130_fd_sc_hs__fill_2 FILLER_49_380 ();
 sky130_fd_sc_hs__fill_1 FILLER_49_382 ();
 sky130_fd_sc_hs__fill_4 FILLER_49_401 ();
 sky130_fd_sc_hs__fill_1 FILLER_49_405 ();
 sky130_fd_sc_hs__fill_4 FILLER_49_407 ();
 sky130_fd_sc_hs__fill_1 FILLER_49_411 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_430 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_438 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_446 ();
 sky130_fd_sc_hs__fill_4 FILLER_49_454 ();
 sky130_fd_sc_hs__fill_2 FILLER_49_458 ();
 sky130_fd_sc_hs__fill_1 FILLER_49_460 ();
 sky130_fd_sc_hs__fill_2 FILLER_49_465 ();
 sky130_fd_sc_hs__fill_1 FILLER_49_467 ();
 sky130_fd_sc_hs__fill_4 FILLER_49_478 ();
 sky130_fd_sc_hs__fill_1 FILLER_49_482 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_509 ();
 sky130_fd_sc_hs__fill_4 FILLER_49_517 ();
 sky130_fd_sc_hs__fill_1 FILLER_49_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_49_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_49_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_50_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_50_28 ();
 sky130_fd_sc_hs__fill_1 FILLER_50_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_39 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_47 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_55 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_63 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_71 ();
 sky130_fd_sc_hs__fill_4 FILLER_50_79 ();
 sky130_fd_sc_hs__fill_1 FILLER_50_86 ();
 sky130_fd_sc_hs__fill_4 FILLER_50_109 ();
 sky130_fd_sc_hs__fill_2 FILLER_50_113 ();
 sky130_fd_sc_hs__fill_2 FILLER_50_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_50_138 ();
 sky130_fd_sc_hs__fill_4 FILLER_50_146 ();
 sky130_fd_sc_hs__fill_1 FILLER_50_150 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_154 ();
 sky130_fd_sc_hs__fill_4 FILLER_50_162 ();
 sky130_fd_sc_hs__fill_2 FILLER_50_166 ();
 sky130_fd_sc_hs__fill_4 FILLER_50_171 ();
 sky130_fd_sc_hs__fill_4 FILLER_50_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_204 ();
 sky130_fd_sc_hs__fill_4 FILLER_50_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_243 ();
 sky130_fd_sc_hs__fill_2 FILLER_50_251 ();
 sky130_fd_sc_hs__fill_1 FILLER_50_253 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_270 ();
 sky130_fd_sc_hs__fill_2 FILLER_50_278 ();
 sky130_fd_sc_hs__fill_2 FILLER_50_316 ();
 sky130_fd_sc_hs__fill_1 FILLER_50_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_328 ();
 sky130_fd_sc_hs__fill_4 FILLER_50_336 ();
 sky130_fd_sc_hs__fill_1 FILLER_50_340 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_359 ();
 sky130_fd_sc_hs__fill_2 FILLER_50_367 ();
 sky130_fd_sc_hs__fill_4 FILLER_50_372 ();
 sky130_fd_sc_hs__fill_1 FILLER_50_376 ();
 sky130_fd_sc_hs__fill_4 FILLER_50_378 ();
 sky130_fd_sc_hs__fill_1 FILLER_50_382 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_419 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_427 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_444 ();
 sky130_fd_sc_hs__fill_4 FILLER_50_452 ();
 sky130_fd_sc_hs__fill_2 FILLER_50_456 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_479 ();
 sky130_fd_sc_hs__fill_4 FILLER_50_487 ();
 sky130_fd_sc_hs__fill_2 FILLER_50_491 ();
 sky130_fd_sc_hs__fill_4 FILLER_50_494 ();
 sky130_fd_sc_hs__fill_2 FILLER_50_498 ();
 sky130_fd_sc_hs__fill_2 FILLER_50_503 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_508 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_516 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_524 ();
 sky130_fd_sc_hs__fill_8 FILLER_50_532 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_16 ();
 sky130_fd_sc_hs__fill_2 FILLER_51_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_51_26 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_35 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_43 ();
 sky130_fd_sc_hs__fill_4 FILLER_51_51 ();
 sky130_fd_sc_hs__fill_2 FILLER_51_55 ();
 sky130_fd_sc_hs__fill_1 FILLER_51_57 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_75 ();
 sky130_fd_sc_hs__fill_4 FILLER_51_83 ();
 sky130_fd_sc_hs__fill_2 FILLER_51_87 ();
 sky130_fd_sc_hs__fill_1 FILLER_51_89 ();
 sky130_fd_sc_hs__fill_4 FILLER_51_108 ();
 sky130_fd_sc_hs__fill_1 FILLER_51_112 ();
 sky130_fd_sc_hs__fill_1 FILLER_51_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_124 ();
 sky130_fd_sc_hs__fill_4 FILLER_51_132 ();
 sky130_fd_sc_hs__fill_2 FILLER_51_136 ();
 sky130_fd_sc_hs__fill_4 FILLER_51_141 ();
 sky130_fd_sc_hs__fill_1 FILLER_51_145 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_51_173 ();
 sky130_fd_sc_hs__fill_4 FILLER_51_175 ();
 sky130_fd_sc_hs__fill_1 FILLER_51_179 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_191 ();
 sky130_fd_sc_hs__fill_2 FILLER_51_199 ();
 sky130_fd_sc_hs__fill_4 FILLER_51_227 ();
 sky130_fd_sc_hs__fill_1 FILLER_51_231 ();
 sky130_fd_sc_hs__fill_1 FILLER_51_233 ();
 sky130_fd_sc_hs__fill_2 FILLER_51_239 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_246 ();
 sky130_fd_sc_hs__fill_1 FILLER_51_254 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_51_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_51_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_357 ();
 sky130_fd_sc_hs__fill_2 FILLER_51_365 ();
 sky130_fd_sc_hs__fill_1 FILLER_51_367 ();
 sky130_fd_sc_hs__fill_2 FILLER_51_404 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_488 ();
 sky130_fd_sc_hs__fill_8 FILLER_51_496 ();
 sky130_fd_sc_hs__fill_4 FILLER_51_504 ();
 sky130_fd_sc_hs__fill_2 FILLER_51_508 ();
 sky130_fd_sc_hs__fill_4 FILLER_51_518 ();
 sky130_fd_sc_hs__fill_2 FILLER_51_523 ();
 sky130_fd_sc_hs__fill_1 FILLER_51_525 ();
 sky130_fd_sc_hs__fill_4 FILLER_51_534 ();
 sky130_fd_sc_hs__fill_2 FILLER_51_538 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_8 ();
 sky130_fd_sc_hs__fill_4 FILLER_52_16 ();
 sky130_fd_sc_hs__fill_1 FILLER_52_20 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_64 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_72 ();
 sky130_fd_sc_hs__fill_4 FILLER_52_80 ();
 sky130_fd_sc_hs__fill_2 FILLER_52_84 ();
 sky130_fd_sc_hs__fill_1 FILLER_52_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_88 ();
 sky130_fd_sc_hs__fill_1 FILLER_52_96 ();
 sky130_fd_sc_hs__fill_4 FILLER_52_100 ();
 sky130_fd_sc_hs__fill_2 FILLER_52_104 ();
 sky130_fd_sc_hs__fill_4 FILLER_52_127 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_134 ();
 sky130_fd_sc_hs__fill_2 FILLER_52_142 ();
 sky130_fd_sc_hs__fill_1 FILLER_52_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_154 ();
 sky130_fd_sc_hs__fill_4 FILLER_52_162 ();
 sky130_fd_sc_hs__fill_1 FILLER_52_166 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_185 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_193 ();
 sky130_fd_sc_hs__fill_2 FILLER_52_201 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_220 ();
 sky130_fd_sc_hs__fill_1 FILLER_52_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_234 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_242 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_250 ();
 sky130_fd_sc_hs__fill_2 FILLER_52_258 ();
 sky130_fd_sc_hs__fill_1 FILLER_52_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_262 ();
 sky130_fd_sc_hs__fill_1 FILLER_52_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_297 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_305 ();
 sky130_fd_sc_hs__fill_4 FILLER_52_313 ();
 sky130_fd_sc_hs__fill_2 FILLER_52_317 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_328 ();
 sky130_fd_sc_hs__fill_4 FILLER_52_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_343 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_351 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_378 ();
 sky130_fd_sc_hs__fill_1 FILLER_52_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_390 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_398 ();
 sky130_fd_sc_hs__fill_4 FILLER_52_409 ();
 sky130_fd_sc_hs__fill_1 FILLER_52_413 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_481 ();
 sky130_fd_sc_hs__fill_4 FILLER_52_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_52_526 ();
 sky130_fd_sc_hs__fill_4 FILLER_52_534 ();
 sky130_fd_sc_hs__fill_2 FILLER_52_538 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_53_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_59 ();
 sky130_fd_sc_hs__fill_4 FILLER_53_67 ();
 sky130_fd_sc_hs__fill_2 FILLER_53_71 ();
 sky130_fd_sc_hs__fill_1 FILLER_53_73 ();
 sky130_fd_sc_hs__fill_4 FILLER_53_77 ();
 sky130_fd_sc_hs__fill_1 FILLER_53_84 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_88 ();
 sky130_fd_sc_hs__fill_4 FILLER_53_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_103 ();
 sky130_fd_sc_hs__fill_4 FILLER_53_111 ();
 sky130_fd_sc_hs__fill_1 FILLER_53_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_53_173 ();
 sky130_fd_sc_hs__fill_4 FILLER_53_175 ();
 sky130_fd_sc_hs__fill_2 FILLER_53_179 ();
 sky130_fd_sc_hs__fill_1 FILLER_53_181 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_193 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_201 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_209 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_217 ();
 sky130_fd_sc_hs__fill_4 FILLER_53_225 ();
 sky130_fd_sc_hs__fill_2 FILLER_53_229 ();
 sky130_fd_sc_hs__fill_1 FILLER_53_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_236 ();
 sky130_fd_sc_hs__fill_1 FILLER_53_244 ();
 sky130_fd_sc_hs__fill_4 FILLER_53_248 ();
 sky130_fd_sc_hs__fill_1 FILLER_53_252 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_256 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_264 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_272 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_280 ();
 sky130_fd_sc_hs__fill_2 FILLER_53_288 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_291 ();
 sky130_fd_sc_hs__fill_4 FILLER_53_299 ();
 sky130_fd_sc_hs__fill_2 FILLER_53_303 ();
 sky130_fd_sc_hs__fill_4 FILLER_53_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_53_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_439 ();
 sky130_fd_sc_hs__fill_2 FILLER_53_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_452 ();
 sky130_fd_sc_hs__fill_4 FILLER_53_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_489 ();
 sky130_fd_sc_hs__fill_1 FILLER_53_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_53_503 ();
 sky130_fd_sc_hs__fill_2 FILLER_53_511 ();
 sky130_fd_sc_hs__fill_1 FILLER_53_521 ();
 sky130_fd_sc_hs__fill_4 FILLER_53_523 ();
 sky130_fd_sc_hs__fill_2 FILLER_53_527 ();
 sky130_fd_sc_hs__fill_1 FILLER_53_529 ();
 sky130_fd_sc_hs__fill_2 FILLER_53_538 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_54_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_54_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_30 ();
 sky130_fd_sc_hs__fill_4 FILLER_54_38 ();
 sky130_fd_sc_hs__fill_1 FILLER_54_42 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_61 ();
 sky130_fd_sc_hs__fill_2 FILLER_54_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_93 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_101 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_109 ();
 sky130_fd_sc_hs__fill_2 FILLER_54_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_125 ();
 sky130_fd_sc_hs__fill_2 FILLER_54_133 ();
 sky130_fd_sc_hs__fill_4 FILLER_54_138 ();
 sky130_fd_sc_hs__fill_2 FILLER_54_142 ();
 sky130_fd_sc_hs__fill_1 FILLER_54_144 ();
 sky130_fd_sc_hs__fill_1 FILLER_54_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_168 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_176 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_184 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_192 ();
 sky130_fd_sc_hs__fill_2 FILLER_54_200 ();
 sky130_fd_sc_hs__fill_1 FILLER_54_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_204 ();
 sky130_fd_sc_hs__fill_2 FILLER_54_212 ();
 sky130_fd_sc_hs__fill_4 FILLER_54_225 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_232 ();
 sky130_fd_sc_hs__fill_4 FILLER_54_240 ();
 sky130_fd_sc_hs__fill_4 FILLER_54_262 ();
 sky130_fd_sc_hs__fill_2 FILLER_54_266 ();
 sky130_fd_sc_hs__fill_1 FILLER_54_268 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_272 ();
 sky130_fd_sc_hs__fill_1 FILLER_54_280 ();
 sky130_fd_sc_hs__fill_4 FILLER_54_287 ();
 sky130_fd_sc_hs__fill_2 FILLER_54_291 ();
 sky130_fd_sc_hs__fill_1 FILLER_54_293 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_297 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_305 ();
 sky130_fd_sc_hs__fill_2 FILLER_54_313 ();
 sky130_fd_sc_hs__fill_1 FILLER_54_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_328 ();
 sky130_fd_sc_hs__fill_1 FILLER_54_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_340 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_348 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_356 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_364 ();
 sky130_fd_sc_hs__fill_4 FILLER_54_372 ();
 sky130_fd_sc_hs__fill_1 FILLER_54_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_417 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_425 ();
 sky130_fd_sc_hs__fill_2 FILLER_54_433 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_436 ();
 sky130_fd_sc_hs__fill_1 FILLER_54_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_448 ();
 sky130_fd_sc_hs__fill_8 FILLER_54_456 ();
 sky130_fd_sc_hs__fill_4 FILLER_54_464 ();
 sky130_fd_sc_hs__fill_2 FILLER_54_468 ();
 sky130_fd_sc_hs__fill_2 FILLER_54_503 ();
 sky130_fd_sc_hs__fill_1 FILLER_54_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_0 ();
 sky130_fd_sc_hs__fill_4 FILLER_55_8 ();
 sky130_fd_sc_hs__fill_2 FILLER_55_12 ();
 sky130_fd_sc_hs__fill_1 FILLER_55_14 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_31 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_39 ();
 sky130_fd_sc_hs__fill_4 FILLER_55_47 ();
 sky130_fd_sc_hs__fill_4 FILLER_55_54 ();
 sky130_fd_sc_hs__fill_4 FILLER_55_59 ();
 sky130_fd_sc_hs__fill_2 FILLER_55_63 ();
 sky130_fd_sc_hs__fill_1 FILLER_55_65 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_90 ();
 sky130_fd_sc_hs__fill_4 FILLER_55_98 ();
 sky130_fd_sc_hs__fill_1 FILLER_55_102 ();
 sky130_fd_sc_hs__fill_4 FILLER_55_109 ();
 sky130_fd_sc_hs__fill_2 FILLER_55_113 ();
 sky130_fd_sc_hs__fill_1 FILLER_55_115 ();
 sky130_fd_sc_hs__fill_1 FILLER_55_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_139 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_147 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_155 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_163 ();
 sky130_fd_sc_hs__fill_2 FILLER_55_171 ();
 sky130_fd_sc_hs__fill_1 FILLER_55_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_191 ();
 sky130_fd_sc_hs__fill_4 FILLER_55_199 ();
 sky130_fd_sc_hs__fill_2 FILLER_55_203 ();
 sky130_fd_sc_hs__fill_1 FILLER_55_205 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_217 ();
 sky130_fd_sc_hs__fill_2 FILLER_55_225 ();
 sky130_fd_sc_hs__fill_2 FILLER_55_230 ();
 sky130_fd_sc_hs__fill_4 FILLER_55_291 ();
 sky130_fd_sc_hs__fill_1 FILLER_55_298 ();
 sky130_fd_sc_hs__fill_2 FILLER_55_317 ();
 sky130_fd_sc_hs__fill_2 FILLER_55_340 ();
 sky130_fd_sc_hs__fill_2 FILLER_55_345 ();
 sky130_fd_sc_hs__fill_1 FILLER_55_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_367 ();
 sky130_fd_sc_hs__fill_4 FILLER_55_375 ();
 sky130_fd_sc_hs__fill_2 FILLER_55_379 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_387 ();
 sky130_fd_sc_hs__fill_4 FILLER_55_395 ();
 sky130_fd_sc_hs__fill_2 FILLER_55_399 ();
 sky130_fd_sc_hs__fill_2 FILLER_55_404 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_425 ();
 sky130_fd_sc_hs__fill_1 FILLER_55_433 ();
 sky130_fd_sc_hs__fill_8 FILLER_55_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_55_463 ();
 sky130_fd_sc_hs__fill_2 FILLER_55_483 ();
 sky130_fd_sc_hs__fill_1 FILLER_55_485 ();
 sky130_fd_sc_hs__fill_2 FILLER_55_500 ();
 sky130_fd_sc_hs__fill_1 FILLER_55_502 ();
 sky130_fd_sc_hs__fill_1 FILLER_55_521 ();
 sky130_fd_sc_hs__fill_4 FILLER_55_533 ();
 sky130_fd_sc_hs__fill_2 FILLER_55_537 ();
 sky130_fd_sc_hs__fill_1 FILLER_55_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_56_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_56_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_46 ();
 sky130_fd_sc_hs__fill_1 FILLER_56_54 ();
 sky130_fd_sc_hs__fill_1 FILLER_56_76 ();
 sky130_fd_sc_hs__fill_4 FILLER_56_83 ();
 sky130_fd_sc_hs__fill_2 FILLER_56_88 ();
 sky130_fd_sc_hs__fill_2 FILLER_56_96 ();
 sky130_fd_sc_hs__fill_1 FILLER_56_98 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_120 ();
 sky130_fd_sc_hs__fill_2 FILLER_56_128 ();
 sky130_fd_sc_hs__fill_4 FILLER_56_140 ();
 sky130_fd_sc_hs__fill_1 FILLER_56_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_162 ();
 sky130_fd_sc_hs__fill_4 FILLER_56_170 ();
 sky130_fd_sc_hs__fill_2 FILLER_56_174 ();
 sky130_fd_sc_hs__fill_4 FILLER_56_187 ();
 sky130_fd_sc_hs__fill_2 FILLER_56_191 ();
 sky130_fd_sc_hs__fill_1 FILLER_56_193 ();
 sky130_fd_sc_hs__fill_4 FILLER_56_197 ();
 sky130_fd_sc_hs__fill_2 FILLER_56_201 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_56_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_262 ();
 sky130_fd_sc_hs__fill_4 FILLER_56_270 ();
 sky130_fd_sc_hs__fill_2 FILLER_56_274 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_279 ();
 sky130_fd_sc_hs__fill_4 FILLER_56_287 ();
 sky130_fd_sc_hs__fill_2 FILLER_56_291 ();
 sky130_fd_sc_hs__fill_1 FILLER_56_293 ();
 sky130_fd_sc_hs__fill_2 FILLER_56_306 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_311 ();
 sky130_fd_sc_hs__fill_4 FILLER_56_320 ();
 sky130_fd_sc_hs__fill_1 FILLER_56_324 ();
 sky130_fd_sc_hs__fill_4 FILLER_56_328 ();
 sky130_fd_sc_hs__fill_2 FILLER_56_332 ();
 sky130_fd_sc_hs__fill_1 FILLER_56_334 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_338 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_365 ();
 sky130_fd_sc_hs__fill_4 FILLER_56_373 ();
 sky130_fd_sc_hs__fill_4 FILLER_56_378 ();
 sky130_fd_sc_hs__fill_2 FILLER_56_382 ();
 sky130_fd_sc_hs__fill_1 FILLER_56_387 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_391 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_399 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_56_434 ();
 sky130_fd_sc_hs__fill_4 FILLER_56_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_458 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_466 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_474 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_482 ();
 sky130_fd_sc_hs__fill_2 FILLER_56_490 ();
 sky130_fd_sc_hs__fill_1 FILLER_56_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_494 ();
 sky130_fd_sc_hs__fill_2 FILLER_56_502 ();
 sky130_fd_sc_hs__fill_1 FILLER_56_504 ();
 sky130_fd_sc_hs__fill_8 FILLER_56_508 ();
 sky130_fd_sc_hs__fill_1 FILLER_56_516 ();
 sky130_fd_sc_hs__fill_4 FILLER_56_535 ();
 sky130_fd_sc_hs__fill_1 FILLER_56_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_59 ();
 sky130_fd_sc_hs__fill_1 FILLER_57_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_71 ();
 sky130_fd_sc_hs__fill_2 FILLER_57_82 ();
 sky130_fd_sc_hs__fill_1 FILLER_57_84 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_106 ();
 sky130_fd_sc_hs__fill_2 FILLER_57_114 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_125 ();
 sky130_fd_sc_hs__fill_4 FILLER_57_133 ();
 sky130_fd_sc_hs__fill_2 FILLER_57_137 ();
 sky130_fd_sc_hs__fill_1 FILLER_57_139 ();
 sky130_fd_sc_hs__fill_4 FILLER_57_161 ();
 sky130_fd_sc_hs__fill_1 FILLER_57_165 ();
 sky130_fd_sc_hs__fill_4 FILLER_57_169 ();
 sky130_fd_sc_hs__fill_1 FILLER_57_173 ();
 sky130_fd_sc_hs__fill_1 FILLER_57_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_179 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_187 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_195 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_224 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_233 ();
 sky130_fd_sc_hs__fill_2 FILLER_57_241 ();
 sky130_fd_sc_hs__fill_1 FILLER_57_243 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_57_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_307 ();
 sky130_fd_sc_hs__fill_4 FILLER_57_315 ();
 sky130_fd_sc_hs__fill_1 FILLER_57_319 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_332 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_340 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_360 ();
 sky130_fd_sc_hs__fill_2 FILLER_57_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_57_370 ();
 sky130_fd_sc_hs__fill_4 FILLER_57_374 ();
 sky130_fd_sc_hs__fill_2 FILLER_57_378 ();
 sky130_fd_sc_hs__fill_2 FILLER_57_383 ();
 sky130_fd_sc_hs__fill_2 FILLER_57_403 ();
 sky130_fd_sc_hs__fill_1 FILLER_57_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_407 ();
 sky130_fd_sc_hs__fill_2 FILLER_57_415 ();
 sky130_fd_sc_hs__fill_1 FILLER_57_417 ();
 sky130_fd_sc_hs__fill_2 FILLER_57_421 ();
 sky130_fd_sc_hs__fill_1 FILLER_57_423 ();
 sky130_fd_sc_hs__fill_4 FILLER_57_442 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_465 ();
 sky130_fd_sc_hs__fill_4 FILLER_57_473 ();
 sky130_fd_sc_hs__fill_2 FILLER_57_477 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_482 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_498 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_506 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_57_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_57_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_8 ();
 sky130_fd_sc_hs__fill_4 FILLER_58_16 ();
 sky130_fd_sc_hs__fill_1 FILLER_58_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_58_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_88 ();
 sky130_fd_sc_hs__fill_4 FILLER_58_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_105 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_113 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_121 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_129 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_137 ();
 sky130_fd_sc_hs__fill_2 FILLER_58_146 ();
 sky130_fd_sc_hs__fill_1 FILLER_58_148 ();
 sky130_fd_sc_hs__fill_1 FILLER_58_156 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_176 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_184 ();
 sky130_fd_sc_hs__fill_2 FILLER_58_192 ();
 sky130_fd_sc_hs__fill_4 FILLER_58_197 ();
 sky130_fd_sc_hs__fill_2 FILLER_58_201 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_215 ();
 sky130_fd_sc_hs__fill_4 FILLER_58_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_58_227 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_240 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_248 ();
 sky130_fd_sc_hs__fill_4 FILLER_58_256 ();
 sky130_fd_sc_hs__fill_1 FILLER_58_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_262 ();
 sky130_fd_sc_hs__fill_4 FILLER_58_270 ();
 sky130_fd_sc_hs__fill_2 FILLER_58_274 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_288 ();
 sky130_fd_sc_hs__fill_4 FILLER_58_296 ();
 sky130_fd_sc_hs__fill_2 FILLER_58_300 ();
 sky130_fd_sc_hs__fill_1 FILLER_58_302 ();
 sky130_fd_sc_hs__fill_4 FILLER_58_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_58_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_386 ();
 sky130_fd_sc_hs__fill_4 FILLER_58_394 ();
 sky130_fd_sc_hs__fill_2 FILLER_58_401 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_421 ();
 sky130_fd_sc_hs__fill_4 FILLER_58_429 ();
 sky130_fd_sc_hs__fill_2 FILLER_58_433 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_58_492 ();
 sky130_fd_sc_hs__fill_4 FILLER_58_515 ();
 sky130_fd_sc_hs__fill_1 FILLER_58_519 ();
 sky130_fd_sc_hs__fill_8 FILLER_58_527 ();
 sky130_fd_sc_hs__fill_4 FILLER_58_535 ();
 sky130_fd_sc_hs__fill_1 FILLER_58_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_32 ();
 sky130_fd_sc_hs__fill_2 FILLER_59_40 ();
 sky130_fd_sc_hs__fill_1 FILLER_59_42 ();
 sky130_fd_sc_hs__fill_2 FILLER_59_46 ();
 sky130_fd_sc_hs__fill_1 FILLER_59_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_63 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_71 ();
 sky130_fd_sc_hs__fill_1 FILLER_59_79 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_59_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_141 ();
 sky130_fd_sc_hs__fill_2 FILLER_59_149 ();
 sky130_fd_sc_hs__fill_1 FILLER_59_151 ();
 sky130_fd_sc_hs__fill_4 FILLER_59_175 ();
 sky130_fd_sc_hs__fill_2 FILLER_59_179 ();
 sky130_fd_sc_hs__fill_1 FILLER_59_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_220 ();
 sky130_fd_sc_hs__fill_4 FILLER_59_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_233 ();
 sky130_fd_sc_hs__fill_1 FILLER_59_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_59_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_59_347 ();
 sky130_fd_sc_hs__fill_4 FILLER_59_349 ();
 sky130_fd_sc_hs__fill_4 FILLER_59_368 ();
 sky130_fd_sc_hs__fill_2 FILLER_59_372 ();
 sky130_fd_sc_hs__fill_1 FILLER_59_374 ();
 sky130_fd_sc_hs__fill_4 FILLER_59_399 ();
 sky130_fd_sc_hs__fill_2 FILLER_59_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_412 ();
 sky130_fd_sc_hs__fill_4 FILLER_59_420 ();
 sky130_fd_sc_hs__fill_2 FILLER_59_424 ();
 sky130_fd_sc_hs__fill_1 FILLER_59_426 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_430 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_438 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_446 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_454 ();
 sky130_fd_sc_hs__fill_2 FILLER_59_462 ();
 sky130_fd_sc_hs__fill_2 FILLER_59_465 ();
 sky130_fd_sc_hs__fill_1 FILLER_59_467 ();
 sky130_fd_sc_hs__fill_2 FILLER_59_520 ();
 sky130_fd_sc_hs__fill_8 FILLER_59_523 ();
 sky130_fd_sc_hs__fill_1 FILLER_59_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_8 ();
 sky130_fd_sc_hs__fill_1 FILLER_60_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_60_25 ();
 sky130_fd_sc_hs__fill_4 FILLER_60_30 ();
 sky130_fd_sc_hs__fill_2 FILLER_60_34 ();
 sky130_fd_sc_hs__fill_4 FILLER_60_72 ();
 sky130_fd_sc_hs__fill_2 FILLER_60_76 ();
 sky130_fd_sc_hs__fill_1 FILLER_60_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_92 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_100 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_108 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_116 ();
 sky130_fd_sc_hs__fill_4 FILLER_60_124 ();
 sky130_fd_sc_hs__fill_2 FILLER_60_128 ();
 sky130_fd_sc_hs__fill_2 FILLER_60_142 ();
 sky130_fd_sc_hs__fill_1 FILLER_60_144 ();
 sky130_fd_sc_hs__fill_2 FILLER_60_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_60_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_228 ();
 sky130_fd_sc_hs__fill_1 FILLER_60_236 ();
 sky130_fd_sc_hs__fill_4 FILLER_60_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_306 ();
 sky130_fd_sc_hs__fill_4 FILLER_60_314 ();
 sky130_fd_sc_hs__fill_1 FILLER_60_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_60_376 ();
 sky130_fd_sc_hs__fill_1 FILLER_60_378 ();
 sky130_fd_sc_hs__fill_4 FILLER_60_397 ();
 sky130_fd_sc_hs__fill_2 FILLER_60_401 ();
 sky130_fd_sc_hs__fill_4 FILLER_60_406 ();
 sky130_fd_sc_hs__fill_4 FILLER_60_428 ();
 sky130_fd_sc_hs__fill_2 FILLER_60_432 ();
 sky130_fd_sc_hs__fill_1 FILLER_60_434 ();
 sky130_fd_sc_hs__fill_4 FILLER_60_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_476 ();
 sky130_fd_sc_hs__fill_4 FILLER_60_484 ();
 sky130_fd_sc_hs__fill_2 FILLER_60_488 ();
 sky130_fd_sc_hs__fill_8 FILLER_60_494 ();
 sky130_fd_sc_hs__fill_4 FILLER_60_502 ();
 sky130_fd_sc_hs__fill_1 FILLER_60_506 ();
 sky130_fd_sc_hs__fill_4 FILLER_60_528 ();
 sky130_fd_sc_hs__fill_4 FILLER_61_0 ();
 sky130_fd_sc_hs__fill_2 FILLER_61_4 ();
 sky130_fd_sc_hs__fill_1 FILLER_61_6 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_15 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_23 ();
 sky130_fd_sc_hs__fill_4 FILLER_61_31 ();
 sky130_fd_sc_hs__fill_2 FILLER_61_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_105 ();
 sky130_fd_sc_hs__fill_2 FILLER_61_113 ();
 sky130_fd_sc_hs__fill_1 FILLER_61_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_125 ();
 sky130_fd_sc_hs__fill_2 FILLER_61_158 ();
 sky130_fd_sc_hs__fill_1 FILLER_61_160 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_199 ();
 sky130_fd_sc_hs__fill_4 FILLER_61_207 ();
 sky130_fd_sc_hs__fill_1 FILLER_61_211 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_61_231 ();
 sky130_fd_sc_hs__fill_4 FILLER_61_233 ();
 sky130_fd_sc_hs__fill_1 FILLER_61_237 ();
 sky130_fd_sc_hs__fill_2 FILLER_61_267 ();
 sky130_fd_sc_hs__fill_1 FILLER_61_269 ();
 sky130_fd_sc_hs__fill_4 FILLER_61_273 ();
 sky130_fd_sc_hs__fill_2 FILLER_61_277 ();
 sky130_fd_sc_hs__fill_2 FILLER_61_304 ();
 sky130_fd_sc_hs__fill_1 FILLER_61_306 ();
 sky130_fd_sc_hs__fill_1 FILLER_61_312 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_326 ();
 sky130_fd_sc_hs__fill_4 FILLER_61_334 ();
 sky130_fd_sc_hs__fill_2 FILLER_61_338 ();
 sky130_fd_sc_hs__fill_1 FILLER_61_340 ();
 sky130_fd_sc_hs__fill_1 FILLER_61_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_357 ();
 sky130_fd_sc_hs__fill_4 FILLER_61_365 ();
 sky130_fd_sc_hs__fill_2 FILLER_61_369 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_61_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_407 ();
 sky130_fd_sc_hs__fill_4 FILLER_61_415 ();
 sky130_fd_sc_hs__fill_1 FILLER_61_419 ();
 sky130_fd_sc_hs__fill_2 FILLER_61_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_61_489 ();
 sky130_fd_sc_hs__fill_2 FILLER_61_497 ();
 sky130_fd_sc_hs__fill_1 FILLER_61_523 ();
 sky130_fd_sc_hs__fill_4 FILLER_61_527 ();
 sky130_fd_sc_hs__fill_1 FILLER_61_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_62_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_62_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_54 ();
 sky130_fd_sc_hs__fill_1 FILLER_62_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_62_144 ();
 sky130_fd_sc_hs__fill_4 FILLER_62_146 ();
 sky130_fd_sc_hs__fill_2 FILLER_62_150 ();
 sky130_fd_sc_hs__fill_1 FILLER_62_152 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_166 ();
 sky130_fd_sc_hs__fill_4 FILLER_62_174 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_62_202 ();
 sky130_fd_sc_hs__fill_4 FILLER_62_204 ();
 sky130_fd_sc_hs__fill_1 FILLER_62_208 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_227 ();
 sky130_fd_sc_hs__fill_2 FILLER_62_235 ();
 sky130_fd_sc_hs__fill_1 FILLER_62_237 ();
 sky130_fd_sc_hs__fill_2 FILLER_62_258 ();
 sky130_fd_sc_hs__fill_1 FILLER_62_260 ();
 sky130_fd_sc_hs__fill_4 FILLER_62_262 ();
 sky130_fd_sc_hs__fill_2 FILLER_62_266 ();
 sky130_fd_sc_hs__fill_4 FILLER_62_297 ();
 sky130_fd_sc_hs__fill_2 FILLER_62_309 ();
 sky130_fd_sc_hs__fill_4 FILLER_62_326 ();
 sky130_fd_sc_hs__fill_2 FILLER_62_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_361 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_369 ();
 sky130_fd_sc_hs__fill_4 FILLER_62_378 ();
 sky130_fd_sc_hs__fill_2 FILLER_62_382 ();
 sky130_fd_sc_hs__fill_1 FILLER_62_384 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_388 ();
 sky130_fd_sc_hs__fill_2 FILLER_62_432 ();
 sky130_fd_sc_hs__fill_1 FILLER_62_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_444 ();
 sky130_fd_sc_hs__fill_2 FILLER_62_452 ();
 sky130_fd_sc_hs__fill_1 FILLER_62_454 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_481 ();
 sky130_fd_sc_hs__fill_4 FILLER_62_489 ();
 sky130_fd_sc_hs__fill_4 FILLER_62_494 ();
 sky130_fd_sc_hs__fill_1 FILLER_62_498 ();
 sky130_fd_sc_hs__fill_8 FILLER_62_502 ();
 sky130_fd_sc_hs__fill_4 FILLER_62_536 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_63_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_76 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_84 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_92 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_100 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_108 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_149 ();
 sky130_fd_sc_hs__fill_2 FILLER_63_157 ();
 sky130_fd_sc_hs__fill_1 FILLER_63_159 ();
 sky130_fd_sc_hs__fill_1 FILLER_63_167 ();
 sky130_fd_sc_hs__fill_2 FILLER_63_171 ();
 sky130_fd_sc_hs__fill_1 FILLER_63_173 ();
 sky130_fd_sc_hs__fill_2 FILLER_63_175 ();
 sky130_fd_sc_hs__fill_4 FILLER_63_195 ();
 sky130_fd_sc_hs__fill_1 FILLER_63_199 ();
 sky130_fd_sc_hs__fill_1 FILLER_63_203 ();
 sky130_fd_sc_hs__fill_2 FILLER_63_229 ();
 sky130_fd_sc_hs__fill_1 FILLER_63_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_241 ();
 sky130_fd_sc_hs__fill_1 FILLER_63_249 ();
 sky130_fd_sc_hs__fill_2 FILLER_63_272 ();
 sky130_fd_sc_hs__fill_1 FILLER_63_274 ();
 sky130_fd_sc_hs__fill_2 FILLER_63_278 ();
 sky130_fd_sc_hs__fill_2 FILLER_63_291 ();
 sky130_fd_sc_hs__fill_1 FILLER_63_293 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_304 ();
 sky130_fd_sc_hs__fill_4 FILLER_63_312 ();
 sky130_fd_sc_hs__fill_2 FILLER_63_316 ();
 sky130_fd_sc_hs__fill_2 FILLER_63_345 ();
 sky130_fd_sc_hs__fill_1 FILLER_63_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_364 ();
 sky130_fd_sc_hs__fill_4 FILLER_63_372 ();
 sky130_fd_sc_hs__fill_1 FILLER_63_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_380 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_423 ();
 sky130_fd_sc_hs__fill_2 FILLER_63_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_452 ();
 sky130_fd_sc_hs__fill_4 FILLER_63_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_473 ();
 sky130_fd_sc_hs__fill_2 FILLER_63_481 ();
 sky130_fd_sc_hs__fill_2 FILLER_63_486 ();
 sky130_fd_sc_hs__fill_1 FILLER_63_488 ();
 sky130_fd_sc_hs__fill_8 FILLER_63_507 ();
 sky130_fd_sc_hs__fill_4 FILLER_63_515 ();
 sky130_fd_sc_hs__fill_2 FILLER_63_519 ();
 sky130_fd_sc_hs__fill_1 FILLER_63_521 ();
 sky130_fd_sc_hs__fill_2 FILLER_63_523 ();
 sky130_fd_sc_hs__fill_2 FILLER_64_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_10 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_18 ();
 sky130_fd_sc_hs__fill_2 FILLER_64_26 ();
 sky130_fd_sc_hs__fill_1 FILLER_64_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_46 ();
 sky130_fd_sc_hs__fill_4 FILLER_64_54 ();
 sky130_fd_sc_hs__fill_1 FILLER_64_58 ();
 sky130_fd_sc_hs__fill_4 FILLER_64_80 ();
 sky130_fd_sc_hs__fill_2 FILLER_64_84 ();
 sky130_fd_sc_hs__fill_1 FILLER_64_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_64_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_154 ();
 sky130_fd_sc_hs__fill_2 FILLER_64_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_181 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_189 ();
 sky130_fd_sc_hs__fill_4 FILLER_64_197 ();
 sky130_fd_sc_hs__fill_2 FILLER_64_201 ();
 sky130_fd_sc_hs__fill_4 FILLER_64_204 ();
 sky130_fd_sc_hs__fill_1 FILLER_64_208 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_249 ();
 sky130_fd_sc_hs__fill_4 FILLER_64_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_262 ();
 sky130_fd_sc_hs__fill_4 FILLER_64_270 ();
 sky130_fd_sc_hs__fill_1 FILLER_64_286 ();
 sky130_fd_sc_hs__fill_4 FILLER_64_295 ();
 sky130_fd_sc_hs__fill_2 FILLER_64_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_307 ();
 sky130_fd_sc_hs__fill_4 FILLER_64_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_344 ();
 sky130_fd_sc_hs__fill_2 FILLER_64_352 ();
 sky130_fd_sc_hs__fill_2 FILLER_64_359 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_369 ();
 sky130_fd_sc_hs__fill_1 FILLER_64_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_382 ();
 sky130_fd_sc_hs__fill_2 FILLER_64_390 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_404 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_412 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_420 ();
 sky130_fd_sc_hs__fill_4 FILLER_64_428 ();
 sky130_fd_sc_hs__fill_2 FILLER_64_432 ();
 sky130_fd_sc_hs__fill_1 FILLER_64_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_64_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_64_510 ();
 sky130_fd_sc_hs__fill_4 FILLER_64_518 ();
 sky130_fd_sc_hs__fill_2 FILLER_64_522 ();
 sky130_fd_sc_hs__fill_1 FILLER_64_524 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_65_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_59 ();
 sky130_fd_sc_hs__fill_2 FILLER_65_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_77 ();
 sky130_fd_sc_hs__fill_4 FILLER_65_85 ();
 sky130_fd_sc_hs__fill_1 FILLER_65_89 ();
 sky130_fd_sc_hs__fill_1 FILLER_65_100 ();
 sky130_fd_sc_hs__fill_2 FILLER_65_113 ();
 sky130_fd_sc_hs__fill_1 FILLER_65_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_129 ();
 sky130_fd_sc_hs__fill_2 FILLER_65_137 ();
 sky130_fd_sc_hs__fill_1 FILLER_65_168 ();
 sky130_fd_sc_hs__fill_1 FILLER_65_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_194 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_252 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_268 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_276 ();
 sky130_fd_sc_hs__fill_4 FILLER_65_284 ();
 sky130_fd_sc_hs__fill_2 FILLER_65_288 ();
 sky130_fd_sc_hs__fill_4 FILLER_65_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_301 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_309 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_317 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_325 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_333 ();
 sky130_fd_sc_hs__fill_4 FILLER_65_341 ();
 sky130_fd_sc_hs__fill_2 FILLER_65_345 ();
 sky130_fd_sc_hs__fill_1 FILLER_65_347 ();
 sky130_fd_sc_hs__fill_1 FILLER_65_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_364 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_372 ();
 sky130_fd_sc_hs__fill_1 FILLER_65_380 ();
 sky130_fd_sc_hs__fill_4 FILLER_65_399 ();
 sky130_fd_sc_hs__fill_2 FILLER_65_403 ();
 sky130_fd_sc_hs__fill_1 FILLER_65_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_447 ();
 sky130_fd_sc_hs__fill_2 FILLER_65_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_65_457 ();
 sky130_fd_sc_hs__fill_4 FILLER_65_483 ();
 sky130_fd_sc_hs__fill_1 FILLER_65_487 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_491 ();
 sky130_fd_sc_hs__fill_4 FILLER_65_499 ();
 sky130_fd_sc_hs__fill_2 FILLER_65_506 ();
 sky130_fd_sc_hs__fill_8 FILLER_65_511 ();
 sky130_fd_sc_hs__fill_2 FILLER_65_519 ();
 sky130_fd_sc_hs__fill_1 FILLER_65_521 ();
 sky130_fd_sc_hs__fill_2 FILLER_65_523 ();
 sky130_fd_sc_hs__fill_4 FILLER_65_536 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_66_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_66_28 ();
 sky130_fd_sc_hs__fill_4 FILLER_66_30 ();
 sky130_fd_sc_hs__fill_1 FILLER_66_34 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_56 ();
 sky130_fd_sc_hs__fill_4 FILLER_66_67 ();
 sky130_fd_sc_hs__fill_2 FILLER_66_71 ();
 sky130_fd_sc_hs__fill_1 FILLER_66_86 ();
 sky130_fd_sc_hs__fill_2 FILLER_66_88 ();
 sky130_fd_sc_hs__fill_1 FILLER_66_90 ();
 sky130_fd_sc_hs__fill_4 FILLER_66_94 ();
 sky130_fd_sc_hs__fill_2 FILLER_66_98 ();
 sky130_fd_sc_hs__fill_4 FILLER_66_141 ();
 sky130_fd_sc_hs__fill_1 FILLER_66_146 ();
 sky130_fd_sc_hs__fill_4 FILLER_66_158 ();
 sky130_fd_sc_hs__fill_2 FILLER_66_162 ();
 sky130_fd_sc_hs__fill_1 FILLER_66_164 ();
 sky130_fd_sc_hs__fill_1 FILLER_66_174 ();
 sky130_fd_sc_hs__fill_1 FILLER_66_180 ();
 sky130_fd_sc_hs__fill_4 FILLER_66_199 ();
 sky130_fd_sc_hs__fill_4 FILLER_66_204 ();
 sky130_fd_sc_hs__fill_2 FILLER_66_208 ();
 sky130_fd_sc_hs__fill_1 FILLER_66_210 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_229 ();
 sky130_fd_sc_hs__fill_4 FILLER_66_237 ();
 sky130_fd_sc_hs__fill_2 FILLER_66_241 ();
 sky130_fd_sc_hs__fill_1 FILLER_66_243 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_270 ();
 sky130_fd_sc_hs__fill_4 FILLER_66_278 ();
 sky130_fd_sc_hs__fill_2 FILLER_66_282 ();
 sky130_fd_sc_hs__fill_1 FILLER_66_284 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_288 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_296 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_304 ();
 sky130_fd_sc_hs__fill_4 FILLER_66_312 ();
 sky130_fd_sc_hs__fill_2 FILLER_66_316 ();
 sky130_fd_sc_hs__fill_1 FILLER_66_318 ();
 sky130_fd_sc_hs__fill_4 FILLER_66_320 ();
 sky130_fd_sc_hs__fill_2 FILLER_66_324 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_338 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_346 ();
 sky130_fd_sc_hs__fill_1 FILLER_66_354 ();
 sky130_fd_sc_hs__fill_4 FILLER_66_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_378 ();
 sky130_fd_sc_hs__fill_1 FILLER_66_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_66_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_66_434 ();
 sky130_fd_sc_hs__fill_2 FILLER_66_436 ();
 sky130_fd_sc_hs__fill_1 FILLER_66_438 ();
 sky130_fd_sc_hs__fill_2 FILLER_66_460 ();
 sky130_fd_sc_hs__fill_1 FILLER_66_462 ();
 sky130_fd_sc_hs__fill_2 FILLER_66_466 ();
 sky130_fd_sc_hs__fill_1 FILLER_66_468 ();
 sky130_fd_sc_hs__fill_2 FILLER_66_472 ();
 sky130_fd_sc_hs__fill_1 FILLER_66_474 ();
 sky130_fd_sc_hs__fill_4 FILLER_66_512 ();
 sky130_fd_sc_hs__fill_2 FILLER_66_516 ();
 sky130_fd_sc_hs__fill_1 FILLER_66_518 ();
 sky130_fd_sc_hs__fill_4 FILLER_66_526 ();
 sky130_fd_sc_hs__fill_2 FILLER_66_530 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_8 ();
 sky130_fd_sc_hs__fill_4 FILLER_67_16 ();
 sky130_fd_sc_hs__fill_2 FILLER_67_20 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_59 ();
 sky130_fd_sc_hs__fill_2 FILLER_67_67 ();
 sky130_fd_sc_hs__fill_1 FILLER_67_69 ();
 sky130_fd_sc_hs__fill_4 FILLER_67_73 ();
 sky130_fd_sc_hs__fill_2 FILLER_67_77 ();
 sky130_fd_sc_hs__fill_2 FILLER_67_82 ();
 sky130_fd_sc_hs__fill_1 FILLER_67_84 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_103 ();
 sky130_fd_sc_hs__fill_4 FILLER_67_111 ();
 sky130_fd_sc_hs__fill_1 FILLER_67_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_117 ();
 sky130_fd_sc_hs__fill_2 FILLER_67_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_142 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_150 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_158 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_166 ();
 sky130_fd_sc_hs__fill_4 FILLER_67_175 ();
 sky130_fd_sc_hs__fill_1 FILLER_67_179 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_67_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_67_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_291 ();
 sky130_fd_sc_hs__fill_4 FILLER_67_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_310 ();
 sky130_fd_sc_hs__fill_4 FILLER_67_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_335 ();
 sky130_fd_sc_hs__fill_4 FILLER_67_343 ();
 sky130_fd_sc_hs__fill_1 FILLER_67_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_349 ();
 sky130_fd_sc_hs__fill_4 FILLER_67_357 ();
 sky130_fd_sc_hs__fill_2 FILLER_67_361 ();
 sky130_fd_sc_hs__fill_1 FILLER_67_363 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_371 ();
 sky130_fd_sc_hs__fill_1 FILLER_67_405 ();
 sky130_fd_sc_hs__fill_2 FILLER_67_407 ();
 sky130_fd_sc_hs__fill_1 FILLER_67_409 ();
 sky130_fd_sc_hs__fill_1 FILLER_67_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_448 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_456 ();
 sky130_fd_sc_hs__fill_8 FILLER_67_465 ();
 sky130_fd_sc_hs__fill_4 FILLER_67_473 ();
 sky130_fd_sc_hs__fill_2 FILLER_67_477 ();
 sky130_fd_sc_hs__fill_1 FILLER_67_479 ();
 sky130_fd_sc_hs__fill_2 FILLER_67_519 ();
 sky130_fd_sc_hs__fill_1 FILLER_67_521 ();
 sky130_fd_sc_hs__fill_2 FILLER_67_530 ();
 sky130_fd_sc_hs__fill_4 FILLER_68_0 ();
 sky130_fd_sc_hs__fill_2 FILLER_68_4 ();
 sky130_fd_sc_hs__fill_1 FILLER_68_6 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_15 ();
 sky130_fd_sc_hs__fill_4 FILLER_68_23 ();
 sky130_fd_sc_hs__fill_2 FILLER_68_27 ();
 sky130_fd_sc_hs__fill_4 FILLER_68_30 ();
 sky130_fd_sc_hs__fill_2 FILLER_68_34 ();
 sky130_fd_sc_hs__fill_1 FILLER_68_36 ();
 sky130_fd_sc_hs__fill_4 FILLER_68_40 ();
 sky130_fd_sc_hs__fill_2 FILLER_68_44 ();
 sky130_fd_sc_hs__fill_4 FILLER_68_82 ();
 sky130_fd_sc_hs__fill_1 FILLER_68_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_120 ();
 sky130_fd_sc_hs__fill_4 FILLER_68_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_165 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_181 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_189 ();
 sky130_fd_sc_hs__fill_4 FILLER_68_197 ();
 sky130_fd_sc_hs__fill_2 FILLER_68_201 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_68_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_286 ();
 sky130_fd_sc_hs__fill_4 FILLER_68_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_311 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_327 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_335 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_343 ();
 sky130_fd_sc_hs__fill_4 FILLER_68_351 ();
 sky130_fd_sc_hs__fill_2 FILLER_68_355 ();
 sky130_fd_sc_hs__fill_1 FILLER_68_357 ();
 sky130_fd_sc_hs__fill_4 FILLER_68_378 ();
 sky130_fd_sc_hs__fill_1 FILLER_68_382 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_390 ();
 sky130_fd_sc_hs__fill_4 FILLER_68_398 ();
 sky130_fd_sc_hs__fill_1 FILLER_68_402 ();
 sky130_fd_sc_hs__fill_4 FILLER_68_429 ();
 sky130_fd_sc_hs__fill_2 FILLER_68_433 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_460 ();
 sky130_fd_sc_hs__fill_1 FILLER_68_468 ();
 sky130_fd_sc_hs__fill_1 FILLER_68_487 ();
 sky130_fd_sc_hs__fill_2 FILLER_68_491 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_68_502 ();
 sky130_fd_sc_hs__fill_4 FILLER_68_510 ();
 sky130_fd_sc_hs__fill_2 FILLER_68_514 ();
 sky130_fd_sc_hs__fill_1 FILLER_68_516 ();
 sky130_fd_sc_hs__fill_1 FILLER_68_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_40 ();
 sky130_fd_sc_hs__fill_4 FILLER_69_48 ();
 sky130_fd_sc_hs__fill_1 FILLER_69_52 ();
 sky130_fd_sc_hs__fill_2 FILLER_69_56 ();
 sky130_fd_sc_hs__fill_1 FILLER_69_59 ();
 sky130_fd_sc_hs__fill_2 FILLER_69_63 ();
 sky130_fd_sc_hs__fill_1 FILLER_69_65 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_69 ();
 sky130_fd_sc_hs__fill_2 FILLER_69_77 ();
 sky130_fd_sc_hs__fill_1 FILLER_69_79 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_69_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_117 ();
 sky130_fd_sc_hs__fill_4 FILLER_69_125 ();
 sky130_fd_sc_hs__fill_1 FILLER_69_129 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_157 ();
 sky130_fd_sc_hs__fill_2 FILLER_69_165 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_69_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_270 ();
 sky130_fd_sc_hs__fill_4 FILLER_69_278 ();
 sky130_fd_sc_hs__fill_1 FILLER_69_282 ();
 sky130_fd_sc_hs__fill_2 FILLER_69_291 ();
 sky130_fd_sc_hs__fill_1 FILLER_69_293 ();
 sky130_fd_sc_hs__fill_4 FILLER_69_311 ();
 sky130_fd_sc_hs__fill_4 FILLER_69_330 ();
 sky130_fd_sc_hs__fill_2 FILLER_69_334 ();
 sky130_fd_sc_hs__fill_4 FILLER_69_343 ();
 sky130_fd_sc_hs__fill_1 FILLER_69_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_69_405 ();
 sky130_fd_sc_hs__fill_2 FILLER_69_407 ();
 sky130_fd_sc_hs__fill_4 FILLER_69_428 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_450 ();
 sky130_fd_sc_hs__fill_4 FILLER_69_458 ();
 sky130_fd_sc_hs__fill_2 FILLER_69_462 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_489 ();
 sky130_fd_sc_hs__fill_4 FILLER_69_497 ();
 sky130_fd_sc_hs__fill_2 FILLER_69_501 ();
 sky130_fd_sc_hs__fill_1 FILLER_69_521 ();
 sky130_fd_sc_hs__fill_1 FILLER_69_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_69_532 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_70_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_70_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_38 ();
 sky130_fd_sc_hs__fill_2 FILLER_70_46 ();
 sky130_fd_sc_hs__fill_4 FILLER_70_51 ();
 sky130_fd_sc_hs__fill_1 FILLER_70_55 ();
 sky130_fd_sc_hs__fill_1 FILLER_70_77 ();
 sky130_fd_sc_hs__fill_4 FILLER_70_81 ();
 sky130_fd_sc_hs__fill_2 FILLER_70_85 ();
 sky130_fd_sc_hs__fill_4 FILLER_70_88 ();
 sky130_fd_sc_hs__fill_1 FILLER_70_92 ();
 sky130_fd_sc_hs__fill_2 FILLER_70_99 ();
 sky130_fd_sc_hs__fill_1 FILLER_70_101 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_105 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_113 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_121 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_129 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_137 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_70_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_204 ();
 sky130_fd_sc_hs__fill_4 FILLER_70_212 ();
 sky130_fd_sc_hs__fill_2 FILLER_70_221 ();
 sky130_fd_sc_hs__fill_1 FILLER_70_223 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_229 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_237 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_267 ();
 sky130_fd_sc_hs__fill_2 FILLER_70_275 ();
 sky130_fd_sc_hs__fill_2 FILLER_70_282 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_311 ();
 sky130_fd_sc_hs__fill_2 FILLER_70_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_70_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_378 ();
 sky130_fd_sc_hs__fill_1 FILLER_70_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_394 ();
 sky130_fd_sc_hs__fill_2 FILLER_70_402 ();
 sky130_fd_sc_hs__fill_1 FILLER_70_404 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_423 ();
 sky130_fd_sc_hs__fill_4 FILLER_70_431 ();
 sky130_fd_sc_hs__fill_4 FILLER_70_436 ();
 sky130_fd_sc_hs__fill_2 FILLER_70_440 ();
 sky130_fd_sc_hs__fill_1 FILLER_70_442 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_483 ();
 sky130_fd_sc_hs__fill_2 FILLER_70_491 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_502 ();
 sky130_fd_sc_hs__fill_4 FILLER_70_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_70_532 ();
 sky130_fd_sc_hs__fill_4 FILLER_71_0 ();
 sky130_fd_sc_hs__fill_2 FILLER_71_4 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_14 ();
 sky130_fd_sc_hs__fill_4 FILLER_71_30 ();
 sky130_fd_sc_hs__fill_2 FILLER_71_34 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_67 ();
 sky130_fd_sc_hs__fill_4 FILLER_71_75 ();
 sky130_fd_sc_hs__fill_1 FILLER_71_79 ();
 sky130_fd_sc_hs__fill_2 FILLER_71_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_108 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_133 ();
 sky130_fd_sc_hs__fill_2 FILLER_71_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_71_173 ();
 sky130_fd_sc_hs__fill_2 FILLER_71_175 ();
 sky130_fd_sc_hs__fill_1 FILLER_71_177 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_189 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_197 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_205 ();
 sky130_fd_sc_hs__fill_1 FILLER_71_213 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_233 ();
 sky130_fd_sc_hs__fill_4 FILLER_71_251 ();
 sky130_fd_sc_hs__fill_2 FILLER_71_255 ();
 sky130_fd_sc_hs__fill_1 FILLER_71_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_278 ();
 sky130_fd_sc_hs__fill_1 FILLER_71_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_291 ();
 sky130_fd_sc_hs__fill_1 FILLER_71_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_312 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_336 ();
 sky130_fd_sc_hs__fill_4 FILLER_71_344 ();
 sky130_fd_sc_hs__fill_2 FILLER_71_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_368 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_384 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_392 ();
 sky130_fd_sc_hs__fill_4 FILLER_71_400 ();
 sky130_fd_sc_hs__fill_2 FILLER_71_404 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_71_463 ();
 sky130_fd_sc_hs__fill_4 FILLER_71_465 ();
 sky130_fd_sc_hs__fill_2 FILLER_71_469 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_474 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_482 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_490 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_498 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_506 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_71_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_71_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_0 ();
 sky130_fd_sc_hs__fill_1 FILLER_72_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_17 ();
 sky130_fd_sc_hs__fill_4 FILLER_72_25 ();
 sky130_fd_sc_hs__fill_4 FILLER_72_30 ();
 sky130_fd_sc_hs__fill_2 FILLER_72_34 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_54 ();
 sky130_fd_sc_hs__fill_4 FILLER_72_62 ();
 sky130_fd_sc_hs__fill_2 FILLER_72_66 ();
 sky130_fd_sc_hs__fill_1 FILLER_72_68 ();
 sky130_fd_sc_hs__fill_2 FILLER_72_72 ();
 sky130_fd_sc_hs__fill_1 FILLER_72_74 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_72_86 ();
 sky130_fd_sc_hs__fill_2 FILLER_72_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_93 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_101 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_109 ();
 sky130_fd_sc_hs__fill_4 FILLER_72_117 ();
 sky130_fd_sc_hs__fill_2 FILLER_72_121 ();
 sky130_fd_sc_hs__fill_1 FILLER_72_123 ();
 sky130_fd_sc_hs__fill_4 FILLER_72_127 ();
 sky130_fd_sc_hs__fill_2 FILLER_72_131 ();
 sky130_fd_sc_hs__fill_2 FILLER_72_138 ();
 sky130_fd_sc_hs__fill_1 FILLER_72_140 ();
 sky130_fd_sc_hs__fill_1 FILLER_72_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_170 ();
 sky130_fd_sc_hs__fill_4 FILLER_72_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_185 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_193 ();
 sky130_fd_sc_hs__fill_2 FILLER_72_201 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_204 ();
 sky130_fd_sc_hs__fill_2 FILLER_72_212 ();
 sky130_fd_sc_hs__fill_1 FILLER_72_214 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_221 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_229 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_237 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_245 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_253 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_262 ();
 sky130_fd_sc_hs__fill_4 FILLER_72_270 ();
 sky130_fd_sc_hs__fill_2 FILLER_72_274 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_305 ();
 sky130_fd_sc_hs__fill_4 FILLER_72_313 ();
 sky130_fd_sc_hs__fill_2 FILLER_72_317 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_340 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_348 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_356 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_364 ();
 sky130_fd_sc_hs__fill_4 FILLER_72_372 ();
 sky130_fd_sc_hs__fill_1 FILLER_72_376 ();
 sky130_fd_sc_hs__fill_2 FILLER_72_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_400 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_408 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_416 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_424 ();
 sky130_fd_sc_hs__fill_2 FILLER_72_432 ();
 sky130_fd_sc_hs__fill_1 FILLER_72_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_460 ();
 sky130_fd_sc_hs__fill_1 FILLER_72_468 ();
 sky130_fd_sc_hs__fill_4 FILLER_72_487 ();
 sky130_fd_sc_hs__fill_2 FILLER_72_491 ();
 sky130_fd_sc_hs__fill_8 FILLER_72_494 ();
 sky130_fd_sc_hs__fill_1 FILLER_72_502 ();
 sky130_fd_sc_hs__fill_2 FILLER_72_530 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_0 ();
 sky130_fd_sc_hs__fill_4 FILLER_73_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_20 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_36 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_44 ();
 sky130_fd_sc_hs__fill_4 FILLER_73_52 ();
 sky130_fd_sc_hs__fill_2 FILLER_73_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_59 ();
 sky130_fd_sc_hs__fill_1 FILLER_73_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_71 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_79 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_87 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_95 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_103 ();
 sky130_fd_sc_hs__fill_4 FILLER_73_111 ();
 sky130_fd_sc_hs__fill_1 FILLER_73_115 ();
 sky130_fd_sc_hs__fill_2 FILLER_73_117 ();
 sky130_fd_sc_hs__fill_1 FILLER_73_119 ();
 sky130_fd_sc_hs__fill_4 FILLER_73_151 ();
 sky130_fd_sc_hs__fill_1 FILLER_73_155 ();
 sky130_fd_sc_hs__fill_4 FILLER_73_159 ();
 sky130_fd_sc_hs__fill_1 FILLER_73_163 ();
 sky130_fd_sc_hs__fill_2 FILLER_73_193 ();
 sky130_fd_sc_hs__fill_1 FILLER_73_195 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_201 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_209 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_217 ();
 sky130_fd_sc_hs__fill_4 FILLER_73_225 ();
 sky130_fd_sc_hs__fill_2 FILLER_73_229 ();
 sky130_fd_sc_hs__fill_1 FILLER_73_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_254 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_278 ();
 sky130_fd_sc_hs__fill_4 FILLER_73_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_73_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_359 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_367 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_375 ();
 sky130_fd_sc_hs__fill_2 FILLER_73_383 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_423 ();
 sky130_fd_sc_hs__fill_4 FILLER_73_431 ();
 sky130_fd_sc_hs__fill_2 FILLER_73_435 ();
 sky130_fd_sc_hs__fill_1 FILLER_73_437 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_483 ();
 sky130_fd_sc_hs__fill_8 FILLER_73_509 ();
 sky130_fd_sc_hs__fill_4 FILLER_73_517 ();
 sky130_fd_sc_hs__fill_1 FILLER_73_521 ();
 sky130_fd_sc_hs__fill_2 FILLER_73_537 ();
 sky130_fd_sc_hs__fill_1 FILLER_73_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_74_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_74_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_54 ();
 sky130_fd_sc_hs__fill_1 FILLER_74_62 ();
 sky130_fd_sc_hs__fill_4 FILLER_74_81 ();
 sky130_fd_sc_hs__fill_2 FILLER_74_85 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_88 ();
 sky130_fd_sc_hs__fill_4 FILLER_74_104 ();
 sky130_fd_sc_hs__fill_1 FILLER_74_108 ();
 sky130_fd_sc_hs__fill_2 FILLER_74_114 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_119 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_127 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_135 ();
 sky130_fd_sc_hs__fill_2 FILLER_74_143 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_164 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_172 ();
 sky130_fd_sc_hs__fill_2 FILLER_74_225 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_248 ();
 sky130_fd_sc_hs__fill_4 FILLER_74_256 ();
 sky130_fd_sc_hs__fill_1 FILLER_74_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_302 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_310 ();
 sky130_fd_sc_hs__fill_1 FILLER_74_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_344 ();
 sky130_fd_sc_hs__fill_4 FILLER_74_352 ();
 sky130_fd_sc_hs__fill_1 FILLER_74_356 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_378 ();
 sky130_fd_sc_hs__fill_2 FILLER_74_386 ();
 sky130_fd_sc_hs__fill_1 FILLER_74_388 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_402 ();
 sky130_fd_sc_hs__fill_1 FILLER_74_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_424 ();
 sky130_fd_sc_hs__fill_2 FILLER_74_432 ();
 sky130_fd_sc_hs__fill_1 FILLER_74_434 ();
 sky130_fd_sc_hs__fill_2 FILLER_74_436 ();
 sky130_fd_sc_hs__fill_1 FILLER_74_438 ();
 sky130_fd_sc_hs__fill_8 FILLER_74_467 ();
 sky130_fd_sc_hs__fill_2 FILLER_74_494 ();
 sky130_fd_sc_hs__fill_1 FILLER_74_496 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_8 ();
 sky130_fd_sc_hs__fill_4 FILLER_75_16 ();
 sky130_fd_sc_hs__fill_1 FILLER_75_20 ();
 sky130_fd_sc_hs__fill_4 FILLER_75_29 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_45 ();
 sky130_fd_sc_hs__fill_4 FILLER_75_53 ();
 sky130_fd_sc_hs__fill_1 FILLER_75_57 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_59 ();
 sky130_fd_sc_hs__fill_4 FILLER_75_67 ();
 sky130_fd_sc_hs__fill_1 FILLER_75_92 ();
 sky130_fd_sc_hs__fill_2 FILLER_75_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_117 ();
 sky130_fd_sc_hs__fill_2 FILLER_75_125 ();
 sky130_fd_sc_hs__fill_1 FILLER_75_127 ();
 sky130_fd_sc_hs__fill_4 FILLER_75_136 ();
 sky130_fd_sc_hs__fill_2 FILLER_75_140 ();
 sky130_fd_sc_hs__fill_1 FILLER_75_142 ();
 sky130_fd_sc_hs__fill_2 FILLER_75_151 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_156 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_164 ();
 sky130_fd_sc_hs__fill_2 FILLER_75_172 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_199 ();
 sky130_fd_sc_hs__fill_4 FILLER_75_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_219 ();
 sky130_fd_sc_hs__fill_4 FILLER_75_227 ();
 sky130_fd_sc_hs__fill_1 FILLER_75_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_241 ();
 sky130_fd_sc_hs__fill_1 FILLER_75_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_261 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_269 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_280 ();
 sky130_fd_sc_hs__fill_2 FILLER_75_288 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_304 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_312 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_340 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_381 ();
 sky130_fd_sc_hs__fill_4 FILLER_75_389 ();
 sky130_fd_sc_hs__fill_1 FILLER_75_393 ();
 sky130_fd_sc_hs__fill_4 FILLER_75_407 ();
 sky130_fd_sc_hs__fill_1 FILLER_75_411 ();
 sky130_fd_sc_hs__fill_4 FILLER_75_458 ();
 sky130_fd_sc_hs__fill_2 FILLER_75_462 ();
 sky130_fd_sc_hs__fill_2 FILLER_75_465 ();
 sky130_fd_sc_hs__fill_1 FILLER_75_467 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_75_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_75_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_8 ();
 sky130_fd_sc_hs__fill_1 FILLER_76_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_76_25 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_38 ();
 sky130_fd_sc_hs__fill_2 FILLER_76_46 ();
 sky130_fd_sc_hs__fill_1 FILLER_76_66 ();
 sky130_fd_sc_hs__fill_2 FILLER_76_85 ();
 sky130_fd_sc_hs__fill_1 FILLER_76_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_117 ();
 sky130_fd_sc_hs__fill_4 FILLER_76_125 ();
 sky130_fd_sc_hs__fill_1 FILLER_76_129 ();
 sky130_fd_sc_hs__fill_2 FILLER_76_137 ();
 sky130_fd_sc_hs__fill_1 FILLER_76_139 ();
 sky130_fd_sc_hs__fill_2 FILLER_76_143 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_191 ();
 sky130_fd_sc_hs__fill_4 FILLER_76_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_220 ();
 sky130_fd_sc_hs__fill_1 FILLER_76_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_237 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_245 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_253 ();
 sky130_fd_sc_hs__fill_2 FILLER_76_262 ();
 sky130_fd_sc_hs__fill_1 FILLER_76_264 ();
 sky130_fd_sc_hs__fill_4 FILLER_76_282 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_301 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_309 ();
 sky130_fd_sc_hs__fill_2 FILLER_76_317 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_76_376 ();
 sky130_fd_sc_hs__fill_2 FILLER_76_378 ();
 sky130_fd_sc_hs__fill_1 FILLER_76_380 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_397 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_413 ();
 sky130_fd_sc_hs__fill_1 FILLER_76_421 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_444 ();
 sky130_fd_sc_hs__fill_4 FILLER_76_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_76_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_76_492 ();
 sky130_fd_sc_hs__fill_4 FILLER_76_494 ();
 sky130_fd_sc_hs__fill_2 FILLER_76_498 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_40 ();
 sky130_fd_sc_hs__fill_2 FILLER_77_48 ();
 sky130_fd_sc_hs__fill_4 FILLER_77_53 ();
 sky130_fd_sc_hs__fill_1 FILLER_77_57 ();
 sky130_fd_sc_hs__fill_4 FILLER_77_59 ();
 sky130_fd_sc_hs__fill_2 FILLER_77_63 ();
 sky130_fd_sc_hs__fill_1 FILLER_77_65 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_69 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_82 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_90 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_98 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_106 ();
 sky130_fd_sc_hs__fill_2 FILLER_77_114 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_117 ();
 sky130_fd_sc_hs__fill_1 FILLER_77_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_159 ();
 sky130_fd_sc_hs__fill_4 FILLER_77_167 ();
 sky130_fd_sc_hs__fill_2 FILLER_77_171 ();
 sky130_fd_sc_hs__fill_1 FILLER_77_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_207 ();
 sky130_fd_sc_hs__fill_4 FILLER_77_215 ();
 sky130_fd_sc_hs__fill_4 FILLER_77_225 ();
 sky130_fd_sc_hs__fill_2 FILLER_77_229 ();
 sky130_fd_sc_hs__fill_1 FILLER_77_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_241 ();
 sky130_fd_sc_hs__fill_4 FILLER_77_249 ();
 sky130_fd_sc_hs__fill_2 FILLER_77_253 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_275 ();
 sky130_fd_sc_hs__fill_4 FILLER_77_283 ();
 sky130_fd_sc_hs__fill_2 FILLER_77_287 ();
 sky130_fd_sc_hs__fill_1 FILLER_77_289 ();
 sky130_fd_sc_hs__fill_1 FILLER_77_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_309 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_317 ();
 sky130_fd_sc_hs__fill_1 FILLER_77_325 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_77_347 ();
 sky130_fd_sc_hs__fill_4 FILLER_77_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_358 ();
 sky130_fd_sc_hs__fill_1 FILLER_77_366 ();
 sky130_fd_sc_hs__fill_1 FILLER_77_379 ();
 sky130_fd_sc_hs__fill_4 FILLER_77_383 ();
 sky130_fd_sc_hs__fill_2 FILLER_77_387 ();
 sky130_fd_sc_hs__fill_1 FILLER_77_389 ();
 sky130_fd_sc_hs__fill_4 FILLER_77_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_77_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_77_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_77_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_77_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_78_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_78_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_30 ();
 sky130_fd_sc_hs__fill_4 FILLER_78_38 ();
 sky130_fd_sc_hs__fill_1 FILLER_78_42 ();
 sky130_fd_sc_hs__fill_4 FILLER_78_61 ();
 sky130_fd_sc_hs__fill_1 FILLER_78_65 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_128 ();
 sky130_fd_sc_hs__fill_2 FILLER_78_136 ();
 sky130_fd_sc_hs__fill_2 FILLER_78_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_78_202 ();
 sky130_fd_sc_hs__fill_4 FILLER_78_224 ();
 sky130_fd_sc_hs__fill_2 FILLER_78_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_247 ();
 sky130_fd_sc_hs__fill_4 FILLER_78_255 ();
 sky130_fd_sc_hs__fill_2 FILLER_78_259 ();
 sky130_fd_sc_hs__fill_2 FILLER_78_279 ();
 sky130_fd_sc_hs__fill_1 FILLER_78_281 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_285 ();
 sky130_fd_sc_hs__fill_4 FILLER_78_302 ();
 sky130_fd_sc_hs__fill_1 FILLER_78_306 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_310 ();
 sky130_fd_sc_hs__fill_1 FILLER_78_318 ();
 sky130_fd_sc_hs__fill_4 FILLER_78_320 ();
 sky130_fd_sc_hs__fill_2 FILLER_78_329 ();
 sky130_fd_sc_hs__fill_4 FILLER_78_334 ();
 sky130_fd_sc_hs__fill_2 FILLER_78_338 ();
 sky130_fd_sc_hs__fill_4 FILLER_78_361 ();
 sky130_fd_sc_hs__fill_1 FILLER_78_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_393 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_401 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_421 ();
 sky130_fd_sc_hs__fill_4 FILLER_78_429 ();
 sky130_fd_sc_hs__fill_2 FILLER_78_433 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_78_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_78_526 ();
 sky130_fd_sc_hs__fill_4 FILLER_78_534 ();
 sky130_fd_sc_hs__fill_2 FILLER_78_538 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_0 ();
 sky130_fd_sc_hs__fill_2 FILLER_79_8 ();
 sky130_fd_sc_hs__fill_1 FILLER_79_10 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_21 ();
 sky130_fd_sc_hs__fill_2 FILLER_79_40 ();
 sky130_fd_sc_hs__fill_4 FILLER_79_52 ();
 sky130_fd_sc_hs__fill_2 FILLER_79_56 ();
 sky130_fd_sc_hs__fill_4 FILLER_79_59 ();
 sky130_fd_sc_hs__fill_2 FILLER_79_63 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_71 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_79 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_87 ();
 sky130_fd_sc_hs__fill_2 FILLER_79_95 ();
 sky130_fd_sc_hs__fill_1 FILLER_79_97 ();
 sky130_fd_sc_hs__fill_2 FILLER_79_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_148 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_156 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_164 ();
 sky130_fd_sc_hs__fill_2 FILLER_79_172 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_199 ();
 sky130_fd_sc_hs__fill_2 FILLER_79_207 ();
 sky130_fd_sc_hs__fill_1 FILLER_79_209 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_250 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_258 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_266 ();
 sky130_fd_sc_hs__fill_4 FILLER_79_274 ();
 sky130_fd_sc_hs__fill_2 FILLER_79_278 ();
 sky130_fd_sc_hs__fill_1 FILLER_79_289 ();
 sky130_fd_sc_hs__fill_2 FILLER_79_291 ();
 sky130_fd_sc_hs__fill_1 FILLER_79_293 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_308 ();
 sky130_fd_sc_hs__fill_4 FILLER_79_316 ();
 sky130_fd_sc_hs__fill_2 FILLER_79_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_79_347 ();
 sky130_fd_sc_hs__fill_4 FILLER_79_349 ();
 sky130_fd_sc_hs__fill_2 FILLER_79_356 ();
 sky130_fd_sc_hs__fill_1 FILLER_79_358 ();
 sky130_fd_sc_hs__fill_4 FILLER_79_374 ();
 sky130_fd_sc_hs__fill_2 FILLER_79_378 ();
 sky130_fd_sc_hs__fill_1 FILLER_79_380 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_394 ();
 sky130_fd_sc_hs__fill_4 FILLER_79_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_407 ();
 sky130_fd_sc_hs__fill_4 FILLER_79_415 ();
 sky130_fd_sc_hs__fill_2 FILLER_79_419 ();
 sky130_fd_sc_hs__fill_1 FILLER_79_421 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_447 ();
 sky130_fd_sc_hs__fill_1 FILLER_79_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_79_463 ();
 sky130_fd_sc_hs__fill_2 FILLER_79_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_478 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_486 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_79_510 ();
 sky130_fd_sc_hs__fill_4 FILLER_79_518 ();
 sky130_fd_sc_hs__fill_4 FILLER_79_523 ();
 sky130_fd_sc_hs__fill_1 FILLER_79_527 ();
 sky130_fd_sc_hs__fill_4 FILLER_79_536 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_8 ();
 sky130_fd_sc_hs__fill_4 FILLER_80_16 ();
 sky130_fd_sc_hs__fill_1 FILLER_80_20 ();
 sky130_fd_sc_hs__fill_1 FILLER_80_48 ();
 sky130_fd_sc_hs__fill_4 FILLER_80_55 ();
 sky130_fd_sc_hs__fill_1 FILLER_80_59 ();
 sky130_fd_sc_hs__fill_4 FILLER_80_78 ();
 sky130_fd_sc_hs__fill_2 FILLER_80_82 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_101 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_109 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_133 ();
 sky130_fd_sc_hs__fill_4 FILLER_80_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_80_202 ();
 sky130_fd_sc_hs__fill_2 FILLER_80_204 ();
 sky130_fd_sc_hs__fill_1 FILLER_80_206 ();
 sky130_fd_sc_hs__fill_4 FILLER_80_256 ();
 sky130_fd_sc_hs__fill_1 FILLER_80_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_270 ();
 sky130_fd_sc_hs__fill_2 FILLER_80_278 ();
 sky130_fd_sc_hs__fill_1 FILLER_80_280 ();
 sky130_fd_sc_hs__fill_4 FILLER_80_284 ();
 sky130_fd_sc_hs__fill_2 FILLER_80_288 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_295 ();
 sky130_fd_sc_hs__fill_4 FILLER_80_303 ();
 sky130_fd_sc_hs__fill_4 FILLER_80_314 ();
 sky130_fd_sc_hs__fill_1 FILLER_80_318 ();
 sky130_fd_sc_hs__fill_1 FILLER_80_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_338 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_346 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_354 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_362 ();
 sky130_fd_sc_hs__fill_4 FILLER_80_370 ();
 sky130_fd_sc_hs__fill_2 FILLER_80_374 ();
 sky130_fd_sc_hs__fill_1 FILLER_80_376 ();
 sky130_fd_sc_hs__fill_4 FILLER_80_378 ();
 sky130_fd_sc_hs__fill_2 FILLER_80_382 ();
 sky130_fd_sc_hs__fill_1 FILLER_80_401 ();
 sky130_fd_sc_hs__fill_2 FILLER_80_411 ();
 sky130_fd_sc_hs__fill_1 FILLER_80_413 ();
 sky130_fd_sc_hs__fill_1 FILLER_80_417 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_424 ();
 sky130_fd_sc_hs__fill_2 FILLER_80_432 ();
 sky130_fd_sc_hs__fill_1 FILLER_80_434 ();
 sky130_fd_sc_hs__fill_4 FILLER_80_436 ();
 sky130_fd_sc_hs__fill_2 FILLER_80_440 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_485 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_80_526 ();
 sky130_fd_sc_hs__fill_4 FILLER_80_534 ();
 sky130_fd_sc_hs__fill_2 FILLER_80_538 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_24 ();
 sky130_fd_sc_hs__fill_4 FILLER_81_32 ();
 sky130_fd_sc_hs__fill_2 FILLER_81_36 ();
 sky130_fd_sc_hs__fill_2 FILLER_81_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_75 ();
 sky130_fd_sc_hs__fill_4 FILLER_81_83 ();
 sky130_fd_sc_hs__fill_1 FILLER_81_87 ();
 sky130_fd_sc_hs__fill_2 FILLER_81_91 ();
 sky130_fd_sc_hs__fill_1 FILLER_81_93 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_97 ();
 sky130_fd_sc_hs__fill_4 FILLER_81_105 ();
 sky130_fd_sc_hs__fill_4 FILLER_81_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_141 ();
 sky130_fd_sc_hs__fill_4 FILLER_81_149 ();
 sky130_fd_sc_hs__fill_1 FILLER_81_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_197 ();
 sky130_fd_sc_hs__fill_4 FILLER_81_205 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_221 ();
 sky130_fd_sc_hs__fill_2 FILLER_81_229 ();
 sky130_fd_sc_hs__fill_1 FILLER_81_231 ();
 sky130_fd_sc_hs__fill_4 FILLER_81_251 ();
 sky130_fd_sc_hs__fill_1 FILLER_81_255 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_303 ();
 sky130_fd_sc_hs__fill_4 FILLER_81_311 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_326 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_334 ();
 sky130_fd_sc_hs__fill_1 FILLER_81_342 ();
 sky130_fd_sc_hs__fill_2 FILLER_81_346 ();
 sky130_fd_sc_hs__fill_4 FILLER_81_349 ();
 sky130_fd_sc_hs__fill_1 FILLER_81_353 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_365 ();
 sky130_fd_sc_hs__fill_1 FILLER_81_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_394 ();
 sky130_fd_sc_hs__fill_4 FILLER_81_402 ();
 sky130_fd_sc_hs__fill_4 FILLER_81_407 ();
 sky130_fd_sc_hs__fill_1 FILLER_81_411 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_491 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_499 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_507 ();
 sky130_fd_sc_hs__fill_4 FILLER_81_515 ();
 sky130_fd_sc_hs__fill_2 FILLER_81_519 ();
 sky130_fd_sc_hs__fill_1 FILLER_81_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_81_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_81_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_82_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_82_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_48 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_64 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_72 ();
 sky130_fd_sc_hs__fill_4 FILLER_82_80 ();
 sky130_fd_sc_hs__fill_2 FILLER_82_84 ();
 sky130_fd_sc_hs__fill_1 FILLER_82_86 ();
 sky130_fd_sc_hs__fill_1 FILLER_82_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_107 ();
 sky130_fd_sc_hs__fill_2 FILLER_82_115 ();
 sky130_fd_sc_hs__fill_1 FILLER_82_117 ();
 sky130_fd_sc_hs__fill_4 FILLER_82_131 ();
 sky130_fd_sc_hs__fill_4 FILLER_82_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_171 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_179 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_187 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_195 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_204 ();
 sky130_fd_sc_hs__fill_4 FILLER_82_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_82_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_280 ();
 sky130_fd_sc_hs__fill_1 FILLER_82_288 ();
 sky130_fd_sc_hs__fill_2 FILLER_82_292 ();
 sky130_fd_sc_hs__fill_1 FILLER_82_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_307 ();
 sky130_fd_sc_hs__fill_4 FILLER_82_315 ();
 sky130_fd_sc_hs__fill_2 FILLER_82_320 ();
 sky130_fd_sc_hs__fill_1 FILLER_82_322 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_329 ();
 sky130_fd_sc_hs__fill_4 FILLER_82_337 ();
 sky130_fd_sc_hs__fill_2 FILLER_82_341 ();
 sky130_fd_sc_hs__fill_1 FILLER_82_343 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_351 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_359 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_367 ();
 sky130_fd_sc_hs__fill_2 FILLER_82_375 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_406 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_414 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_422 ();
 sky130_fd_sc_hs__fill_4 FILLER_82_430 ();
 sky130_fd_sc_hs__fill_1 FILLER_82_434 ();
 sky130_fd_sc_hs__fill_4 FILLER_82_440 ();
 sky130_fd_sc_hs__fill_1 FILLER_82_456 ();
 sky130_fd_sc_hs__fill_4 FILLER_82_466 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_82_502 ();
 sky130_fd_sc_hs__fill_4 FILLER_82_510 ();
 sky130_fd_sc_hs__fill_2 FILLER_82_514 ();
 sky130_fd_sc_hs__fill_1 FILLER_82_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_83_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_83_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_83_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_83_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_83_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_83_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_83_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_83_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_83_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_83_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_83_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_83_83 ();
 sky130_fd_sc_hs__fill_4 FILLER_83_91 ();
 sky130_fd_sc_hs__fill_2 FILLER_83_113 ();
 sky130_fd_sc_hs__fill_1 FILLER_83_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_83_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_83_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_83_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_83_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_83_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_83_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_83_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_83_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_83_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_83_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_83_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_83_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_83_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_83_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_83_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_83_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_83_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_83_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_83_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_83_257 ();
 sky130_fd_sc_hs__fill_4 FILLER_83_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_83_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_83_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_83_307 ();
 sky130_fd_sc_hs__fill_4 FILLER_83_315 ();
 sky130_fd_sc_hs__fill_2 FILLER_83_319 ();
 sky130_fd_sc_hs__fill_1 FILLER_83_321 ();
 sky130_fd_sc_hs__fill_8 FILLER_83_335 ();
 sky130_fd_sc_hs__fill_4 FILLER_83_343 ();
 sky130_fd_sc_hs__fill_1 FILLER_83_347 ();
 sky130_fd_sc_hs__fill_2 FILLER_83_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_83_368 ();
 sky130_fd_sc_hs__fill_8 FILLER_83_376 ();
 sky130_fd_sc_hs__fill_4 FILLER_83_384 ();
 sky130_fd_sc_hs__fill_1 FILLER_83_388 ();
 sky130_fd_sc_hs__fill_4 FILLER_83_407 ();
 sky130_fd_sc_hs__fill_1 FILLER_83_411 ();
 sky130_fd_sc_hs__fill_8 FILLER_83_417 ();
 sky130_fd_sc_hs__fill_8 FILLER_83_425 ();
 sky130_fd_sc_hs__fill_8 FILLER_83_433 ();
 sky130_fd_sc_hs__fill_8 FILLER_83_441 ();
 sky130_fd_sc_hs__fill_2 FILLER_83_449 ();
 sky130_fd_sc_hs__fill_8 FILLER_83_454 ();
 sky130_fd_sc_hs__fill_2 FILLER_83_462 ();
 sky130_fd_sc_hs__fill_8 FILLER_83_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_83_473 ();
 sky130_fd_sc_hs__fill_4 FILLER_83_481 ();
 sky130_fd_sc_hs__fill_2 FILLER_83_485 ();
 sky130_fd_sc_hs__fill_1 FILLER_83_487 ();
 sky130_fd_sc_hs__fill_8 FILLER_83_511 ();
 sky130_fd_sc_hs__fill_2 FILLER_83_519 ();
 sky130_fd_sc_hs__fill_1 FILLER_83_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_83_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_83_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_83_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_84_0 ();
 sky130_fd_sc_hs__fill_2 FILLER_84_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_84_18 ();
 sky130_fd_sc_hs__fill_2 FILLER_84_26 ();
 sky130_fd_sc_hs__fill_1 FILLER_84_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_84_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_84_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_84_46 ();
 sky130_fd_sc_hs__fill_4 FILLER_84_54 ();
 sky130_fd_sc_hs__fill_1 FILLER_84_58 ();
 sky130_fd_sc_hs__fill_4 FILLER_84_77 ();
 sky130_fd_sc_hs__fill_2 FILLER_84_81 ();
 sky130_fd_sc_hs__fill_1 FILLER_84_83 ();
 sky130_fd_sc_hs__fill_1 FILLER_84_106 ();
 sky130_fd_sc_hs__fill_8 FILLER_84_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_84_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_84_146 ();
 sky130_fd_sc_hs__fill_4 FILLER_84_154 ();
 sky130_fd_sc_hs__fill_2 FILLER_84_158 ();
 sky130_fd_sc_hs__fill_8 FILLER_84_172 ();
 sky130_fd_sc_hs__fill_2 FILLER_84_180 ();
 sky130_fd_sc_hs__fill_1 FILLER_84_182 ();
 sky130_fd_sc_hs__fill_8 FILLER_84_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_84_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_84_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_84_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_84_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_84_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_84_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_84_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_84_262 ();
 sky130_fd_sc_hs__fill_1 FILLER_84_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_84_285 ();
 sky130_fd_sc_hs__fill_8 FILLER_84_293 ();
 sky130_fd_sc_hs__fill_8 FILLER_84_304 ();
 sky130_fd_sc_hs__fill_2 FILLER_84_312 ();
 sky130_fd_sc_hs__fill_1 FILLER_84_314 ();
 sky130_fd_sc_hs__fill_1 FILLER_84_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_84_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_84_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_84_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_84_344 ();
 sky130_fd_sc_hs__fill_4 FILLER_84_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_84_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_84_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_84_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_84_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_84_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_84_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_84_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_84_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_84_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_84_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_84_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_84_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_84_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_84_476 ();
 sky130_fd_sc_hs__fill_4 FILLER_84_484 ();
 sky130_fd_sc_hs__fill_2 FILLER_84_488 ();
 sky130_fd_sc_hs__fill_8 FILLER_84_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_84_502 ();
 sky130_fd_sc_hs__fill_2 FILLER_84_510 ();
 sky130_fd_sc_hs__fill_4 FILLER_84_535 ();
 sky130_fd_sc_hs__fill_1 FILLER_84_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_85_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_85_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_85_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_85_24 ();
 sky130_fd_sc_hs__fill_2 FILLER_85_32 ();
 sky130_fd_sc_hs__fill_1 FILLER_85_34 ();
 sky130_fd_sc_hs__fill_2 FILLER_85_38 ();
 sky130_fd_sc_hs__fill_2 FILLER_85_59 ();
 sky130_fd_sc_hs__fill_1 FILLER_85_61 ();
 sky130_fd_sc_hs__fill_8 FILLER_85_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_85_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_85_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_85_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_85_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_85_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_85_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_85_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_85_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_85_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_85_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_85_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_85_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_85_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_85_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_85_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_85_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_85_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_85_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_85_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_85_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_85_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_85_245 ();
 sky130_fd_sc_hs__fill_8 FILLER_85_253 ();
 sky130_fd_sc_hs__fill_8 FILLER_85_261 ();
 sky130_fd_sc_hs__fill_8 FILLER_85_269 ();
 sky130_fd_sc_hs__fill_8 FILLER_85_277 ();
 sky130_fd_sc_hs__fill_4 FILLER_85_285 ();
 sky130_fd_sc_hs__fill_1 FILLER_85_289 ();
 sky130_fd_sc_hs__fill_2 FILLER_85_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_85_296 ();
 sky130_fd_sc_hs__fill_2 FILLER_85_304 ();
 sky130_fd_sc_hs__fill_1 FILLER_85_306 ();
 sky130_fd_sc_hs__fill_8 FILLER_85_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_85_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_85_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_85_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_85_349 ();
 sky130_fd_sc_hs__fill_4 FILLER_85_357 ();
 sky130_fd_sc_hs__fill_1 FILLER_85_361 ();
 sky130_fd_sc_hs__fill_1 FILLER_85_384 ();
 sky130_fd_sc_hs__fill_8 FILLER_85_407 ();
 sky130_fd_sc_hs__fill_4 FILLER_85_415 ();
 sky130_fd_sc_hs__fill_1 FILLER_85_419 ();
 sky130_fd_sc_hs__fill_8 FILLER_85_440 ();
 sky130_fd_sc_hs__fill_8 FILLER_85_448 ();
 sky130_fd_sc_hs__fill_8 FILLER_85_456 ();
 sky130_fd_sc_hs__fill_8 FILLER_85_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_85_473 ();
 sky130_fd_sc_hs__fill_2 FILLER_85_481 ();
 sky130_fd_sc_hs__fill_1 FILLER_85_483 ();
 sky130_fd_sc_hs__fill_1 FILLER_85_514 ();
 sky130_fd_sc_hs__fill_4 FILLER_85_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_85_523 ();
 sky130_fd_sc_hs__fill_1 FILLER_85_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_86_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_86_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_86_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_86_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_86_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_86_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_86_38 ();
 sky130_fd_sc_hs__fill_4 FILLER_86_46 ();
 sky130_fd_sc_hs__fill_2 FILLER_86_50 ();
 sky130_fd_sc_hs__fill_1 FILLER_86_52 ();
 sky130_fd_sc_hs__fill_2 FILLER_86_62 ();
 sky130_fd_sc_hs__fill_1 FILLER_86_64 ();
 sky130_fd_sc_hs__fill_8 FILLER_86_68 ();
 sky130_fd_sc_hs__fill_8 FILLER_86_76 ();
 sky130_fd_sc_hs__fill_2 FILLER_86_84 ();
 sky130_fd_sc_hs__fill_1 FILLER_86_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_86_88 ();
 sky130_fd_sc_hs__fill_2 FILLER_86_96 ();
 sky130_fd_sc_hs__fill_1 FILLER_86_98 ();
 sky130_fd_sc_hs__fill_8 FILLER_86_102 ();
 sky130_fd_sc_hs__fill_8 FILLER_86_110 ();
 sky130_fd_sc_hs__fill_8 FILLER_86_118 ();
 sky130_fd_sc_hs__fill_8 FILLER_86_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_86_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_86_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_86_191 ();
 sky130_fd_sc_hs__fill_4 FILLER_86_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_86_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_86_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_86_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_86_249 ();
 sky130_fd_sc_hs__fill_4 FILLER_86_257 ();
 sky130_fd_sc_hs__fill_4 FILLER_86_262 ();
 sky130_fd_sc_hs__fill_2 FILLER_86_266 ();
 sky130_fd_sc_hs__fill_2 FILLER_86_285 ();
 sky130_fd_sc_hs__fill_1 FILLER_86_287 ();
 sky130_fd_sc_hs__fill_2 FILLER_86_301 ();
 sky130_fd_sc_hs__fill_8 FILLER_86_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_86_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_86_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_86_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_86_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_86_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_86_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_86_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_86_378 ();
 sky130_fd_sc_hs__fill_2 FILLER_86_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_86_422 ();
 sky130_fd_sc_hs__fill_4 FILLER_86_430 ();
 sky130_fd_sc_hs__fill_1 FILLER_86_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_86_436 ();
 sky130_fd_sc_hs__fill_4 FILLER_86_444 ();
 sky130_fd_sc_hs__fill_1 FILLER_86_448 ();
 sky130_fd_sc_hs__fill_8 FILLER_86_472 ();
 sky130_fd_sc_hs__fill_4 FILLER_86_480 ();
 sky130_fd_sc_hs__fill_1 FILLER_86_484 ();
 sky130_fd_sc_hs__fill_4 FILLER_86_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_86_497 ();
 sky130_fd_sc_hs__fill_2 FILLER_86_505 ();
 sky130_fd_sc_hs__fill_1 FILLER_86_507 ();
 sky130_fd_sc_hs__fill_8 FILLER_86_516 ();
 sky130_fd_sc_hs__fill_8 FILLER_86_524 ();
 sky130_fd_sc_hs__fill_8 FILLER_86_532 ();
 sky130_fd_sc_hs__fill_4 FILLER_87_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_87_20 ();
 sky130_fd_sc_hs__fill_8 FILLER_87_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_87_36 ();
 sky130_fd_sc_hs__fill_4 FILLER_87_44 ();
 sky130_fd_sc_hs__fill_8 FILLER_87_81 ();
 sky130_fd_sc_hs__fill_4 FILLER_87_89 ();
 sky130_fd_sc_hs__fill_1 FILLER_87_93 ();
 sky130_fd_sc_hs__fill_8 FILLER_87_104 ();
 sky130_fd_sc_hs__fill_4 FILLER_87_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_87_117 ();
 sky130_fd_sc_hs__fill_2 FILLER_87_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_87_153 ();
 sky130_fd_sc_hs__fill_8 FILLER_87_161 ();
 sky130_fd_sc_hs__fill_4 FILLER_87_169 ();
 sky130_fd_sc_hs__fill_1 FILLER_87_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_87_175 ();
 sky130_fd_sc_hs__fill_4 FILLER_87_183 ();
 sky130_fd_sc_hs__fill_1 FILLER_87_187 ();
 sky130_fd_sc_hs__fill_8 FILLER_87_191 ();
 sky130_fd_sc_hs__fill_2 FILLER_87_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_87_204 ();
 sky130_fd_sc_hs__fill_1 FILLER_87_212 ();
 sky130_fd_sc_hs__fill_2 FILLER_87_220 ();
 sky130_fd_sc_hs__fill_4 FILLER_87_225 ();
 sky130_fd_sc_hs__fill_2 FILLER_87_229 ();
 sky130_fd_sc_hs__fill_1 FILLER_87_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_87_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_87_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_87_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_87_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_87_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_87_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_87_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_87_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_87_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_87_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_87_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_87_315 ();
 sky130_fd_sc_hs__fill_2 FILLER_87_323 ();
 sky130_fd_sc_hs__fill_1 FILLER_87_325 ();
 sky130_fd_sc_hs__fill_8 FILLER_87_338 ();
 sky130_fd_sc_hs__fill_2 FILLER_87_346 ();
 sky130_fd_sc_hs__fill_8 FILLER_87_349 ();
 sky130_fd_sc_hs__fill_4 FILLER_87_357 ();
 sky130_fd_sc_hs__fill_2 FILLER_87_361 ();
 sky130_fd_sc_hs__fill_8 FILLER_87_384 ();
 sky130_fd_sc_hs__fill_8 FILLER_87_392 ();
 sky130_fd_sc_hs__fill_4 FILLER_87_400 ();
 sky130_fd_sc_hs__fill_2 FILLER_87_404 ();
 sky130_fd_sc_hs__fill_8 FILLER_87_407 ();
 sky130_fd_sc_hs__fill_4 FILLER_87_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_87_426 ();
 sky130_fd_sc_hs__fill_2 FILLER_87_434 ();
 sky130_fd_sc_hs__fill_1 FILLER_87_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_87_454 ();
 sky130_fd_sc_hs__fill_2 FILLER_87_462 ();
 sky130_fd_sc_hs__fill_8 FILLER_87_488 ();
 sky130_fd_sc_hs__fill_2 FILLER_87_496 ();
 sky130_fd_sc_hs__fill_1 FILLER_87_498 ();
 sky130_fd_sc_hs__fill_8 FILLER_87_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_87_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_87_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_88_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_88_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_88_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_88_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_88_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_88_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_88_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_88_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_88_54 ();
 sky130_fd_sc_hs__fill_4 FILLER_88_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_88_76 ();
 sky130_fd_sc_hs__fill_2 FILLER_88_84 ();
 sky130_fd_sc_hs__fill_1 FILLER_88_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_88_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_88_96 ();
 sky130_fd_sc_hs__fill_2 FILLER_88_104 ();
 sky130_fd_sc_hs__fill_4 FILLER_88_139 ();
 sky130_fd_sc_hs__fill_2 FILLER_88_143 ();
 sky130_fd_sc_hs__fill_8 FILLER_88_146 ();
 sky130_fd_sc_hs__fill_4 FILLER_88_154 ();
 sky130_fd_sc_hs__fill_4 FILLER_88_228 ();
 sky130_fd_sc_hs__fill_1 FILLER_88_232 ();
 sky130_fd_sc_hs__fill_8 FILLER_88_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_88_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_88_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_88_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_88_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_88_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_88_278 ();
 sky130_fd_sc_hs__fill_2 FILLER_88_286 ();
 sky130_fd_sc_hs__fill_1 FILLER_88_288 ();
 sky130_fd_sc_hs__fill_1 FILLER_88_292 ();
 sky130_fd_sc_hs__fill_2 FILLER_88_317 ();
 sky130_fd_sc_hs__fill_8 FILLER_88_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_88_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_88_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_88_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_88_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_88_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_88_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_88_376 ();
 sky130_fd_sc_hs__fill_1 FILLER_88_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_88_422 ();
 sky130_fd_sc_hs__fill_4 FILLER_88_430 ();
 sky130_fd_sc_hs__fill_1 FILLER_88_434 ();
 sky130_fd_sc_hs__fill_2 FILLER_88_436 ();
 sky130_fd_sc_hs__fill_2 FILLER_88_450 ();
 sky130_fd_sc_hs__fill_1 FILLER_88_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_88_479 ();
 sky130_fd_sc_hs__fill_4 FILLER_88_487 ();
 sky130_fd_sc_hs__fill_2 FILLER_88_491 ();
 sky130_fd_sc_hs__fill_8 FILLER_88_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_88_502 ();
 sky130_fd_sc_hs__fill_1 FILLER_88_514 ();
 sky130_fd_sc_hs__fill_2 FILLER_88_538 ();
 sky130_fd_sc_hs__fill_8 FILLER_89_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_89_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_89_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_89_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_89_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_89_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_89_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_89_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_89_59 ();
 sky130_fd_sc_hs__fill_4 FILLER_89_67 ();
 sky130_fd_sc_hs__fill_1 FILLER_89_92 ();
 sky130_fd_sc_hs__fill_2 FILLER_89_114 ();
 sky130_fd_sc_hs__fill_1 FILLER_89_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_89_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_89_154 ();
 sky130_fd_sc_hs__fill_2 FILLER_89_162 ();
 sky130_fd_sc_hs__fill_1 FILLER_89_164 ();
 sky130_fd_sc_hs__fill_4 FILLER_89_168 ();
 sky130_fd_sc_hs__fill_2 FILLER_89_172 ();
 sky130_fd_sc_hs__fill_4 FILLER_89_212 ();
 sky130_fd_sc_hs__fill_2 FILLER_89_216 ();
 sky130_fd_sc_hs__fill_1 FILLER_89_218 ();
 sky130_fd_sc_hs__fill_2 FILLER_89_229 ();
 sky130_fd_sc_hs__fill_1 FILLER_89_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_89_233 ();
 sky130_fd_sc_hs__fill_4 FILLER_89_241 ();
 sky130_fd_sc_hs__fill_1 FILLER_89_251 ();
 sky130_fd_sc_hs__fill_8 FILLER_89_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_89_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_89_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_89_289 ();
 sky130_fd_sc_hs__fill_4 FILLER_89_302 ();
 sky130_fd_sc_hs__fill_2 FILLER_89_306 ();
 sky130_fd_sc_hs__fill_4 FILLER_89_321 ();
 sky130_fd_sc_hs__fill_2 FILLER_89_325 ();
 sky130_fd_sc_hs__fill_2 FILLER_89_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_89_368 ();
 sky130_fd_sc_hs__fill_8 FILLER_89_376 ();
 sky130_fd_sc_hs__fill_1 FILLER_89_384 ();
 sky130_fd_sc_hs__fill_8 FILLER_89_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_89_415 ();
 sky130_fd_sc_hs__fill_1 FILLER_89_423 ();
 sky130_fd_sc_hs__fill_2 FILLER_89_448 ();
 sky130_fd_sc_hs__fill_4 FILLER_89_454 ();
 sky130_fd_sc_hs__fill_2 FILLER_89_458 ();
 sky130_fd_sc_hs__fill_1 FILLER_89_468 ();
 sky130_fd_sc_hs__fill_1 FILLER_89_472 ();
 sky130_fd_sc_hs__fill_2 FILLER_89_493 ();
 sky130_fd_sc_hs__fill_4 FILLER_89_515 ();
 sky130_fd_sc_hs__fill_2 FILLER_89_519 ();
 sky130_fd_sc_hs__fill_1 FILLER_89_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_89_523 ();
 sky130_fd_sc_hs__fill_1 FILLER_89_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_90_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_90_8 ();
 sky130_fd_sc_hs__fill_4 FILLER_90_16 ();
 sky130_fd_sc_hs__fill_1 FILLER_90_20 ();
 sky130_fd_sc_hs__fill_8 FILLER_90_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_90_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_90_46 ();
 sky130_fd_sc_hs__fill_2 FILLER_90_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_90_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_90_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_90_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_90_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_90_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_90_112 ();
 sky130_fd_sc_hs__fill_4 FILLER_90_120 ();
 sky130_fd_sc_hs__fill_2 FILLER_90_124 ();
 sky130_fd_sc_hs__fill_8 FILLER_90_146 ();
 sky130_fd_sc_hs__fill_2 FILLER_90_154 ();
 sky130_fd_sc_hs__fill_4 FILLER_90_193 ();
 sky130_fd_sc_hs__fill_8 FILLER_90_204 ();
 sky130_fd_sc_hs__fill_4 FILLER_90_232 ();
 sky130_fd_sc_hs__fill_1 FILLER_90_236 ();
 sky130_fd_sc_hs__fill_4 FILLER_90_283 ();
 sky130_fd_sc_hs__fill_2 FILLER_90_299 ();
 sky130_fd_sc_hs__fill_1 FILLER_90_301 ();
 sky130_fd_sc_hs__fill_8 FILLER_90_320 ();
 sky130_fd_sc_hs__fill_2 FILLER_90_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_90_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_90_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_90_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_90_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_90_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_90_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_90_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_90_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_90_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_90_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_90_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_90_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_90_456 ();
 sky130_fd_sc_hs__fill_8 FILLER_90_464 ();
 sky130_fd_sc_hs__fill_8 FILLER_90_472 ();
 sky130_fd_sc_hs__fill_8 FILLER_90_480 ();
 sky130_fd_sc_hs__fill_4 FILLER_90_488 ();
 sky130_fd_sc_hs__fill_1 FILLER_90_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_90_494 ();
 sky130_fd_sc_hs__fill_2 FILLER_90_502 ();
 sky130_fd_sc_hs__fill_1 FILLER_90_504 ();
 sky130_fd_sc_hs__fill_8 FILLER_90_508 ();
 sky130_fd_sc_hs__fill_8 FILLER_90_516 ();
 sky130_fd_sc_hs__fill_4 FILLER_90_524 ();
 sky130_fd_sc_hs__fill_1 FILLER_90_528 ();
 sky130_fd_sc_hs__fill_2 FILLER_90_537 ();
 sky130_fd_sc_hs__fill_1 FILLER_90_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_91_0 ();
 sky130_fd_sc_hs__fill_4 FILLER_91_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_91_20 ();
 sky130_fd_sc_hs__fill_8 FILLER_91_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_91_36 ();
 sky130_fd_sc_hs__fill_8 FILLER_91_44 ();
 sky130_fd_sc_hs__fill_4 FILLER_91_52 ();
 sky130_fd_sc_hs__fill_2 FILLER_91_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_91_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_91_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_91_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_91_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_91_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_91_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_91_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_91_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_91_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_91_125 ();
 sky130_fd_sc_hs__fill_4 FILLER_91_133 ();
 sky130_fd_sc_hs__fill_2 FILLER_91_137 ();
 sky130_fd_sc_hs__fill_1 FILLER_91_139 ();
 sky130_fd_sc_hs__fill_8 FILLER_91_152 ();
 sky130_fd_sc_hs__fill_2 FILLER_91_160 ();
 sky130_fd_sc_hs__fill_1 FILLER_91_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_91_166 ();
 sky130_fd_sc_hs__fill_1 FILLER_91_195 ();
 sky130_fd_sc_hs__fill_8 FILLER_91_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_91_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_91_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_91_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_91_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_91_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_91_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_91_249 ();
 sky130_fd_sc_hs__fill_1 FILLER_91_257 ();
 sky130_fd_sc_hs__fill_1 FILLER_91_261 ();
 sky130_fd_sc_hs__fill_8 FILLER_91_269 ();
 sky130_fd_sc_hs__fill_2 FILLER_91_291 ();
 sky130_fd_sc_hs__fill_1 FILLER_91_293 ();
 sky130_fd_sc_hs__fill_8 FILLER_91_297 ();
 sky130_fd_sc_hs__fill_8 FILLER_91_305 ();
 sky130_fd_sc_hs__fill_1 FILLER_91_313 ();
 sky130_fd_sc_hs__fill_2 FILLER_91_324 ();
 sky130_fd_sc_hs__fill_1 FILLER_91_326 ();
 sky130_fd_sc_hs__fill_8 FILLER_91_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_91_374 ();
 sky130_fd_sc_hs__fill_8 FILLER_91_382 ();
 sky130_fd_sc_hs__fill_8 FILLER_91_390 ();
 sky130_fd_sc_hs__fill_8 FILLER_91_398 ();
 sky130_fd_sc_hs__fill_8 FILLER_91_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_91_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_91_423 ();
 sky130_fd_sc_hs__fill_4 FILLER_91_431 ();
 sky130_fd_sc_hs__fill_2 FILLER_91_435 ();
 sky130_fd_sc_hs__fill_1 FILLER_91_437 ();
 sky130_fd_sc_hs__fill_8 FILLER_91_451 ();
 sky130_fd_sc_hs__fill_4 FILLER_91_459 ();
 sky130_fd_sc_hs__fill_1 FILLER_91_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_91_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_91_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_91_481 ();
 sky130_fd_sc_hs__fill_2 FILLER_91_493 ();
 sky130_fd_sc_hs__fill_4 FILLER_91_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_91_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_91_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_91_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_92_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_92_8 ();
 sky130_fd_sc_hs__fill_4 FILLER_92_16 ();
 sky130_fd_sc_hs__fill_1 FILLER_92_20 ();
 sky130_fd_sc_hs__fill_8 FILLER_92_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_92_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_92_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_92_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_92_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_92_70 ();
 sky130_fd_sc_hs__fill_4 FILLER_92_81 ();
 sky130_fd_sc_hs__fill_2 FILLER_92_85 ();
 sky130_fd_sc_hs__fill_8 FILLER_92_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_92_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_92_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_92_112 ();
 sky130_fd_sc_hs__fill_4 FILLER_92_120 ();
 sky130_fd_sc_hs__fill_2 FILLER_92_124 ();
 sky130_fd_sc_hs__fill_1 FILLER_92_126 ();
 sky130_fd_sc_hs__fill_8 FILLER_92_132 ();
 sky130_fd_sc_hs__fill_4 FILLER_92_140 ();
 sky130_fd_sc_hs__fill_1 FILLER_92_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_92_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_92_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_92_162 ();
 sky130_fd_sc_hs__fill_4 FILLER_92_170 ();
 sky130_fd_sc_hs__fill_4 FILLER_92_187 ();
 sky130_fd_sc_hs__fill_2 FILLER_92_191 ();
 sky130_fd_sc_hs__fill_2 FILLER_92_200 ();
 sky130_fd_sc_hs__fill_1 FILLER_92_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_92_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_92_212 ();
 sky130_fd_sc_hs__fill_2 FILLER_92_220 ();
 sky130_fd_sc_hs__fill_1 FILLER_92_222 ();
 sky130_fd_sc_hs__fill_8 FILLER_92_230 ();
 sky130_fd_sc_hs__fill_8 FILLER_92_238 ();
 sky130_fd_sc_hs__fill_8 FILLER_92_246 ();
 sky130_fd_sc_hs__fill_4 FILLER_92_254 ();
 sky130_fd_sc_hs__fill_2 FILLER_92_258 ();
 sky130_fd_sc_hs__fill_1 FILLER_92_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_92_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_92_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_92_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_92_286 ();
 sky130_fd_sc_hs__fill_1 FILLER_92_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_92_308 ();
 sky130_fd_sc_hs__fill_2 FILLER_92_316 ();
 sky130_fd_sc_hs__fill_1 FILLER_92_318 ();
 sky130_fd_sc_hs__fill_4 FILLER_92_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_92_341 ();
 sky130_fd_sc_hs__fill_8 FILLER_92_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_92_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_92_365 ();
 sky130_fd_sc_hs__fill_4 FILLER_92_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_92_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_92_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_92_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_92_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_92_410 ();
 sky130_fd_sc_hs__fill_4 FILLER_92_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_92_457 ();
 sky130_fd_sc_hs__fill_8 FILLER_92_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_92_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_92_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_92_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_92_494 ();
 sky130_fd_sc_hs__fill_2 FILLER_92_502 ();
 sky130_fd_sc_hs__fill_1 FILLER_92_504 ();
 sky130_fd_sc_hs__fill_8 FILLER_93_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_93_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_93_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_93_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_93_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_93_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_93_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_93_56 ();
 sky130_fd_sc_hs__fill_4 FILLER_93_59 ();
 sky130_fd_sc_hs__fill_2 FILLER_93_63 ();
 sky130_fd_sc_hs__fill_8 FILLER_93_85 ();
 sky130_fd_sc_hs__fill_8 FILLER_93_93 ();
 sky130_fd_sc_hs__fill_8 FILLER_93_101 ();
 sky130_fd_sc_hs__fill_4 FILLER_93_109 ();
 sky130_fd_sc_hs__fill_2 FILLER_93_113 ();
 sky130_fd_sc_hs__fill_1 FILLER_93_115 ();
 sky130_fd_sc_hs__fill_2 FILLER_93_141 ();
 sky130_fd_sc_hs__fill_4 FILLER_93_169 ();
 sky130_fd_sc_hs__fill_1 FILLER_93_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_93_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_93_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_93_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_93_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_93_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_93_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_93_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_93_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_93_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_93_252 ();
 sky130_fd_sc_hs__fill_8 FILLER_93_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_93_268 ();
 sky130_fd_sc_hs__fill_8 FILLER_93_276 ();
 sky130_fd_sc_hs__fill_4 FILLER_93_284 ();
 sky130_fd_sc_hs__fill_2 FILLER_93_288 ();
 sky130_fd_sc_hs__fill_8 FILLER_93_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_93_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_93_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_93_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_93_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_93_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_93_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_93_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_93_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_93_357 ();
 sky130_fd_sc_hs__fill_4 FILLER_93_365 ();
 sky130_fd_sc_hs__fill_2 FILLER_93_369 ();
 sky130_fd_sc_hs__fill_1 FILLER_93_371 ();
 sky130_fd_sc_hs__fill_8 FILLER_93_393 ();
 sky130_fd_sc_hs__fill_4 FILLER_93_401 ();
 sky130_fd_sc_hs__fill_1 FILLER_93_405 ();
 sky130_fd_sc_hs__fill_2 FILLER_93_407 ();
 sky130_fd_sc_hs__fill_1 FILLER_93_409 ();
 sky130_fd_sc_hs__fill_8 FILLER_93_419 ();
 sky130_fd_sc_hs__fill_8 FILLER_93_427 ();
 sky130_fd_sc_hs__fill_8 FILLER_93_435 ();
 sky130_fd_sc_hs__fill_8 FILLER_93_443 ();
 sky130_fd_sc_hs__fill_8 FILLER_93_451 ();
 sky130_fd_sc_hs__fill_1 FILLER_93_459 ();
 sky130_fd_sc_hs__fill_8 FILLER_93_488 ();
 sky130_fd_sc_hs__fill_8 FILLER_93_496 ();
 sky130_fd_sc_hs__fill_8 FILLER_93_504 ();
 sky130_fd_sc_hs__fill_4 FILLER_93_512 ();
 sky130_fd_sc_hs__fill_2 FILLER_93_519 ();
 sky130_fd_sc_hs__fill_1 FILLER_93_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_93_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_93_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_93_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_94_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_94_8 ();
 sky130_fd_sc_hs__fill_4 FILLER_94_16 ();
 sky130_fd_sc_hs__fill_1 FILLER_94_20 ();
 sky130_fd_sc_hs__fill_8 FILLER_94_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_94_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_94_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_94_54 ();
 sky130_fd_sc_hs__fill_4 FILLER_94_62 ();
 sky130_fd_sc_hs__fill_1 FILLER_94_66 ();
 sky130_fd_sc_hs__fill_8 FILLER_94_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_94_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_94_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_94_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_94_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_94_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_94_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_94_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_94_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_94_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_94_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_94_170 ();
 sky130_fd_sc_hs__fill_4 FILLER_94_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_94_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_94_212 ();
 sky130_fd_sc_hs__fill_1 FILLER_94_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_94_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_94_249 ();
 sky130_fd_sc_hs__fill_4 FILLER_94_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_94_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_94_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_94_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_94_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_94_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_94_302 ();
 sky130_fd_sc_hs__fill_8 FILLER_94_310 ();
 sky130_fd_sc_hs__fill_1 FILLER_94_318 ();
 sky130_fd_sc_hs__fill_1 FILLER_94_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_94_338 ();
 sky130_fd_sc_hs__fill_8 FILLER_94_346 ();
 sky130_fd_sc_hs__fill_8 FILLER_94_354 ();
 sky130_fd_sc_hs__fill_8 FILLER_94_362 ();
 sky130_fd_sc_hs__fill_4 FILLER_94_370 ();
 sky130_fd_sc_hs__fill_2 FILLER_94_374 ();
 sky130_fd_sc_hs__fill_1 FILLER_94_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_94_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_94_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_94_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_94_402 ();
 sky130_fd_sc_hs__fill_4 FILLER_94_410 ();
 sky130_fd_sc_hs__fill_1 FILLER_94_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_94_460 ();
 sky130_fd_sc_hs__fill_2 FILLER_94_468 ();
 sky130_fd_sc_hs__fill_1 FILLER_94_470 ();
 sky130_fd_sc_hs__fill_2 FILLER_94_491 ();
 sky130_fd_sc_hs__fill_4 FILLER_94_506 ();
 sky130_fd_sc_hs__fill_2 FILLER_94_510 ();
 sky130_fd_sc_hs__fill_1 FILLER_94_512 ();
 sky130_fd_sc_hs__fill_8 FILLER_95_0 ();
 sky130_fd_sc_hs__fill_4 FILLER_95_16 ();
 sky130_fd_sc_hs__fill_1 FILLER_95_20 ();
 sky130_fd_sc_hs__fill_8 FILLER_95_28 ();
 sky130_fd_sc_hs__fill_2 FILLER_95_36 ();
 sky130_fd_sc_hs__fill_4 FILLER_95_59 ();
 sky130_fd_sc_hs__fill_2 FILLER_95_63 ();
 sky130_fd_sc_hs__fill_8 FILLER_95_77 ();
 sky130_fd_sc_hs__fill_8 FILLER_95_85 ();
 sky130_fd_sc_hs__fill_8 FILLER_95_93 ();
 sky130_fd_sc_hs__fill_8 FILLER_95_101 ();
 sky130_fd_sc_hs__fill_4 FILLER_95_109 ();
 sky130_fd_sc_hs__fill_2 FILLER_95_113 ();
 sky130_fd_sc_hs__fill_1 FILLER_95_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_95_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_95_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_95_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_95_141 ();
 sky130_fd_sc_hs__fill_4 FILLER_95_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_95_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_95_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_95_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_95_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_95_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_95_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_95_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_95_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_95_233 ();
 sky130_fd_sc_hs__fill_2 FILLER_95_241 ();
 sky130_fd_sc_hs__fill_1 FILLER_95_243 ();
 sky130_fd_sc_hs__fill_4 FILLER_95_247 ();
 sky130_fd_sc_hs__fill_8 FILLER_95_267 ();
 sky130_fd_sc_hs__fill_8 FILLER_95_275 ();
 sky130_fd_sc_hs__fill_4 FILLER_95_283 ();
 sky130_fd_sc_hs__fill_2 FILLER_95_287 ();
 sky130_fd_sc_hs__fill_1 FILLER_95_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_95_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_95_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_95_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_95_315 ();
 sky130_fd_sc_hs__fill_4 FILLER_95_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_95_349 ();
 sky130_fd_sc_hs__fill_4 FILLER_95_357 ();
 sky130_fd_sc_hs__fill_2 FILLER_95_361 ();
 sky130_fd_sc_hs__fill_1 FILLER_95_363 ();
 sky130_fd_sc_hs__fill_8 FILLER_95_407 ();
 sky130_fd_sc_hs__fill_4 FILLER_95_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_95_438 ();
 sky130_fd_sc_hs__fill_8 FILLER_95_446 ();
 sky130_fd_sc_hs__fill_2 FILLER_95_454 ();
 sky130_fd_sc_hs__fill_1 FILLER_95_460 ();
 sky130_fd_sc_hs__fill_2 FILLER_95_488 ();
 sky130_fd_sc_hs__fill_1 FILLER_95_490 ();
 sky130_fd_sc_hs__fill_8 FILLER_95_523 ();
 sky130_fd_sc_hs__fill_1 FILLER_95_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_96_0 ();
 sky130_fd_sc_hs__fill_4 FILLER_96_8 ();
 sky130_fd_sc_hs__fill_2 FILLER_96_12 ();
 sky130_fd_sc_hs__fill_4 FILLER_96_22 ();
 sky130_fd_sc_hs__fill_2 FILLER_96_26 ();
 sky130_fd_sc_hs__fill_1 FILLER_96_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_96_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_96_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_96_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_96_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_96_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_96_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_96_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_96_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_96_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_96_96 ();
 sky130_fd_sc_hs__fill_2 FILLER_96_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_96_126 ();
 sky130_fd_sc_hs__fill_8 FILLER_96_134 ();
 sky130_fd_sc_hs__fill_2 FILLER_96_142 ();
 sky130_fd_sc_hs__fill_1 FILLER_96_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_96_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_96_188 ();
 sky130_fd_sc_hs__fill_4 FILLER_96_196 ();
 sky130_fd_sc_hs__fill_2 FILLER_96_200 ();
 sky130_fd_sc_hs__fill_1 FILLER_96_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_96_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_96_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_96_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_96_228 ();
 sky130_fd_sc_hs__fill_1 FILLER_96_236 ();
 sky130_fd_sc_hs__fill_2 FILLER_96_269 ();
 sky130_fd_sc_hs__fill_1 FILLER_96_271 ();
 sky130_fd_sc_hs__fill_8 FILLER_96_289 ();
 sky130_fd_sc_hs__fill_1 FILLER_96_297 ();
 sky130_fd_sc_hs__fill_8 FILLER_96_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_96_328 ();
 sky130_fd_sc_hs__fill_2 FILLER_96_336 ();
 sky130_fd_sc_hs__fill_1 FILLER_96_338 ();
 sky130_fd_sc_hs__fill_8 FILLER_96_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_96_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_96_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_96_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_96_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_96_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_96_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_96_434 ();
 sky130_fd_sc_hs__fill_4 FILLER_96_442 ();
 sky130_fd_sc_hs__fill_2 FILLER_96_446 ();
 sky130_fd_sc_hs__fill_1 FILLER_96_448 ();
 sky130_fd_sc_hs__fill_4 FILLER_96_482 ();
 sky130_fd_sc_hs__fill_2 FILLER_96_486 ();
 sky130_fd_sc_hs__fill_2 FILLER_96_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_96_522 ();
 sky130_fd_sc_hs__fill_8 FILLER_96_530 ();
 sky130_fd_sc_hs__fill_2 FILLER_96_538 ();
 sky130_fd_sc_hs__fill_8 FILLER_97_0 ();
 sky130_fd_sc_hs__fill_4 FILLER_97_8 ();
 sky130_fd_sc_hs__fill_1 FILLER_97_12 ();
 sky130_fd_sc_hs__fill_8 FILLER_97_21 ();
 sky130_fd_sc_hs__fill_8 FILLER_97_29 ();
 sky130_fd_sc_hs__fill_8 FILLER_97_37 ();
 sky130_fd_sc_hs__fill_8 FILLER_97_45 ();
 sky130_fd_sc_hs__fill_4 FILLER_97_53 ();
 sky130_fd_sc_hs__fill_1 FILLER_97_57 ();
 sky130_fd_sc_hs__fill_8 FILLER_97_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_97_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_97_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_97_83 ();
 sky130_fd_sc_hs__fill_4 FILLER_97_91 ();
 sky130_fd_sc_hs__fill_1 FILLER_97_95 ();
 sky130_fd_sc_hs__fill_8 FILLER_97_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_97_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_97_133 ();
 sky130_fd_sc_hs__fill_2 FILLER_97_141 ();
 sky130_fd_sc_hs__fill_4 FILLER_97_155 ();
 sky130_fd_sc_hs__fill_8 FILLER_97_162 ();
 sky130_fd_sc_hs__fill_4 FILLER_97_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_97_175 ();
 sky130_fd_sc_hs__fill_1 FILLER_97_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_97_187 ();
 sky130_fd_sc_hs__fill_1 FILLER_97_195 ();
 sky130_fd_sc_hs__fill_8 FILLER_97_220 ();
 sky130_fd_sc_hs__fill_4 FILLER_97_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_97_233 ();
 sky130_fd_sc_hs__fill_4 FILLER_97_241 ();
 sky130_fd_sc_hs__fill_1 FILLER_97_245 ();
 sky130_fd_sc_hs__fill_8 FILLER_97_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_97_257 ();
 sky130_fd_sc_hs__fill_4 FILLER_97_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_97_333 ();
 sky130_fd_sc_hs__fill_4 FILLER_97_341 ();
 sky130_fd_sc_hs__fill_2 FILLER_97_345 ();
 sky130_fd_sc_hs__fill_1 FILLER_97_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_97_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_97_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_97_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_97_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_97_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_97_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_97_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_97_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_97_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_97_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_97_423 ();
 sky130_fd_sc_hs__fill_4 FILLER_97_431 ();
 sky130_fd_sc_hs__fill_2 FILLER_97_435 ();
 sky130_fd_sc_hs__fill_1 FILLER_97_437 ();
 sky130_fd_sc_hs__fill_2 FILLER_97_461 ();
 sky130_fd_sc_hs__fill_1 FILLER_97_463 ();
 sky130_fd_sc_hs__fill_4 FILLER_97_465 ();
 sky130_fd_sc_hs__fill_1 FILLER_97_469 ();
 sky130_fd_sc_hs__fill_8 FILLER_97_476 ();
 sky130_fd_sc_hs__fill_4 FILLER_97_484 ();
 sky130_fd_sc_hs__fill_4 FILLER_97_515 ();
 sky130_fd_sc_hs__fill_2 FILLER_97_519 ();
 sky130_fd_sc_hs__fill_1 FILLER_97_521 ();
 sky130_fd_sc_hs__fill_1 FILLER_97_523 ();
 sky130_fd_sc_hs__fill_4 FILLER_98_0 ();
 sky130_fd_sc_hs__fill_1 FILLER_98_4 ();
 sky130_fd_sc_hs__fill_8 FILLER_98_13 ();
 sky130_fd_sc_hs__fill_8 FILLER_98_21 ();
 sky130_fd_sc_hs__fill_8 FILLER_98_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_98_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_98_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_98_54 ();
 sky130_fd_sc_hs__fill_4 FILLER_98_62 ();
 sky130_fd_sc_hs__fill_1 FILLER_98_66 ();
 sky130_fd_sc_hs__fill_8 FILLER_98_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_98_96 ();
 sky130_fd_sc_hs__fill_2 FILLER_98_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_98_126 ();
 sky130_fd_sc_hs__fill_8 FILLER_98_134 ();
 sky130_fd_sc_hs__fill_2 FILLER_98_142 ();
 sky130_fd_sc_hs__fill_1 FILLER_98_144 ();
 sky130_fd_sc_hs__fill_4 FILLER_98_146 ();
 sky130_fd_sc_hs__fill_1 FILLER_98_150 ();
 sky130_fd_sc_hs__fill_8 FILLER_98_184 ();
 sky130_fd_sc_hs__fill_8 FILLER_98_192 ();
 sky130_fd_sc_hs__fill_1 FILLER_98_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_98_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_98_239 ();
 sky130_fd_sc_hs__fill_8 FILLER_98_247 ();
 sky130_fd_sc_hs__fill_4 FILLER_98_255 ();
 sky130_fd_sc_hs__fill_2 FILLER_98_259 ();
 sky130_fd_sc_hs__fill_2 FILLER_98_262 ();
 sky130_fd_sc_hs__fill_1 FILLER_98_264 ();
 sky130_fd_sc_hs__fill_8 FILLER_98_272 ();
 sky130_fd_sc_hs__fill_8 FILLER_98_280 ();
 sky130_fd_sc_hs__fill_8 FILLER_98_288 ();
 sky130_fd_sc_hs__fill_8 FILLER_98_296 ();
 sky130_fd_sc_hs__fill_8 FILLER_98_304 ();
 sky130_fd_sc_hs__fill_4 FILLER_98_312 ();
 sky130_fd_sc_hs__fill_2 FILLER_98_316 ();
 sky130_fd_sc_hs__fill_1 FILLER_98_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_98_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_98_328 ();
 sky130_fd_sc_hs__fill_4 FILLER_98_336 ();
 sky130_fd_sc_hs__fill_1 FILLER_98_340 ();
 sky130_fd_sc_hs__fill_2 FILLER_98_374 ();
 sky130_fd_sc_hs__fill_1 FILLER_98_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_98_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_98_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_98_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_98_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_98_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_98_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_98_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_98_434 ();
 sky130_fd_sc_hs__fill_4 FILLER_98_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_98_443 ();
 sky130_fd_sc_hs__fill_8 FILLER_98_451 ();
 sky130_fd_sc_hs__fill_8 FILLER_98_459 ();
 sky130_fd_sc_hs__fill_8 FILLER_98_467 ();
 sky130_fd_sc_hs__fill_8 FILLER_98_475 ();
 sky130_fd_sc_hs__fill_2 FILLER_98_483 ();
 sky130_fd_sc_hs__fill_1 FILLER_98_485 ();
 sky130_fd_sc_hs__fill_2 FILLER_98_490 ();
 sky130_fd_sc_hs__fill_1 FILLER_98_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_98_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_98_505 ();
 sky130_fd_sc_hs__fill_1 FILLER_98_513 ();
 sky130_fd_sc_hs__fill_8 FILLER_99_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_99_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_99_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_99_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_99_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_99_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_99_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_99_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_99_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_99_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_99_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_99_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_99_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_99_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_99_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_99_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_99_117 ();
 sky130_fd_sc_hs__fill_4 FILLER_99_125 ();
 sky130_fd_sc_hs__fill_4 FILLER_99_132 ();
 sky130_fd_sc_hs__fill_1 FILLER_99_136 ();
 sky130_fd_sc_hs__fill_4 FILLER_99_140 ();
 sky130_fd_sc_hs__fill_8 FILLER_99_147 ();
 sky130_fd_sc_hs__fill_8 FILLER_99_155 ();
 sky130_fd_sc_hs__fill_8 FILLER_99_163 ();
 sky130_fd_sc_hs__fill_2 FILLER_99_171 ();
 sky130_fd_sc_hs__fill_1 FILLER_99_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_99_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_99_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_99_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_99_199 ();
 sky130_fd_sc_hs__fill_4 FILLER_99_207 ();
 sky130_fd_sc_hs__fill_2 FILLER_99_217 ();
 sky130_fd_sc_hs__fill_1 FILLER_99_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_99_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_99_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_99_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_99_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_99_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_99_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_99_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_99_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_99_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_99_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_99_315 ();
 sky130_fd_sc_hs__fill_4 FILLER_99_323 ();
 sky130_fd_sc_hs__fill_2 FILLER_99_327 ();
 sky130_fd_sc_hs__fill_2 FILLER_99_346 ();
 sky130_fd_sc_hs__fill_2 FILLER_99_349 ();
 sky130_fd_sc_hs__fill_1 FILLER_99_351 ();
 sky130_fd_sc_hs__fill_8 FILLER_99_364 ();
 sky130_fd_sc_hs__fill_8 FILLER_99_372 ();
 sky130_fd_sc_hs__fill_8 FILLER_99_380 ();
 sky130_fd_sc_hs__fill_8 FILLER_99_388 ();
 sky130_fd_sc_hs__fill_8 FILLER_99_396 ();
 sky130_fd_sc_hs__fill_2 FILLER_99_404 ();
 sky130_fd_sc_hs__fill_8 FILLER_99_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_99_415 ();
 sky130_fd_sc_hs__fill_4 FILLER_99_436 ();
 sky130_fd_sc_hs__fill_1 FILLER_99_440 ();
 sky130_fd_sc_hs__fill_8 FILLER_99_465 ();
 sky130_fd_sc_hs__fill_4 FILLER_99_473 ();
 sky130_fd_sc_hs__fill_2 FILLER_99_477 ();
 sky130_fd_sc_hs__fill_2 FILLER_99_509 ();
 sky130_fd_sc_hs__fill_1 FILLER_99_511 ();
 sky130_fd_sc_hs__fill_4 FILLER_99_516 ();
 sky130_fd_sc_hs__fill_2 FILLER_99_520 ();
 sky130_fd_sc_hs__fill_1 FILLER_99_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_100_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_100_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_100_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_100_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_100_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_100_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_100_46 ();
 sky130_fd_sc_hs__fill_4 FILLER_100_54 ();
 sky130_fd_sc_hs__fill_1 FILLER_100_58 ();
 sky130_fd_sc_hs__fill_8 FILLER_100_68 ();
 sky130_fd_sc_hs__fill_8 FILLER_100_76 ();
 sky130_fd_sc_hs__fill_2 FILLER_100_84 ();
 sky130_fd_sc_hs__fill_1 FILLER_100_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_100_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_100_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_100_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_100_112 ();
 sky130_fd_sc_hs__fill_4 FILLER_100_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_100_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_100_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_100_162 ();
 sky130_fd_sc_hs__fill_1 FILLER_100_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_100_184 ();
 sky130_fd_sc_hs__fill_8 FILLER_100_192 ();
 sky130_fd_sc_hs__fill_2 FILLER_100_200 ();
 sky130_fd_sc_hs__fill_1 FILLER_100_202 ();
 sky130_fd_sc_hs__fill_4 FILLER_100_204 ();
 sky130_fd_sc_hs__fill_2 FILLER_100_208 ();
 sky130_fd_sc_hs__fill_1 FILLER_100_210 ();
 sky130_fd_sc_hs__fill_8 FILLER_100_218 ();
 sky130_fd_sc_hs__fill_8 FILLER_100_226 ();
 sky130_fd_sc_hs__fill_8 FILLER_100_237 ();
 sky130_fd_sc_hs__fill_8 FILLER_100_245 ();
 sky130_fd_sc_hs__fill_8 FILLER_100_253 ();
 sky130_fd_sc_hs__fill_2 FILLER_100_262 ();
 sky130_fd_sc_hs__fill_1 FILLER_100_264 ();
 sky130_fd_sc_hs__fill_8 FILLER_100_276 ();
 sky130_fd_sc_hs__fill_8 FILLER_100_284 ();
 sky130_fd_sc_hs__fill_8 FILLER_100_292 ();
 sky130_fd_sc_hs__fill_2 FILLER_100_300 ();
 sky130_fd_sc_hs__fill_4 FILLER_100_312 ();
 sky130_fd_sc_hs__fill_2 FILLER_100_316 ();
 sky130_fd_sc_hs__fill_1 FILLER_100_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_100_320 ();
 sky130_fd_sc_hs__fill_4 FILLER_100_328 ();
 sky130_fd_sc_hs__fill_2 FILLER_100_332 ();
 sky130_fd_sc_hs__fill_1 FILLER_100_334 ();
 sky130_fd_sc_hs__fill_1 FILLER_100_356 ();
 sky130_fd_sc_hs__fill_8 FILLER_100_378 ();
 sky130_fd_sc_hs__fill_1 FILLER_100_386 ();
 sky130_fd_sc_hs__fill_1 FILLER_100_408 ();
 sky130_fd_sc_hs__fill_2 FILLER_100_430 ();
 sky130_fd_sc_hs__fill_4 FILLER_100_444 ();
 sky130_fd_sc_hs__fill_1 FILLER_100_448 ();
 sky130_fd_sc_hs__fill_8 FILLER_100_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_100_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_100_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_100_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_100_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_100_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_100_494 ();
 sky130_fd_sc_hs__fill_1 FILLER_100_502 ();
 sky130_fd_sc_hs__fill_4 FILLER_100_507 ();
 sky130_fd_sc_hs__fill_2 FILLER_100_511 ();
 sky130_fd_sc_hs__fill_4 FILLER_100_536 ();
 sky130_fd_sc_hs__fill_4 FILLER_101_0 ();
 sky130_fd_sc_hs__fill_1 FILLER_101_4 ();
 sky130_fd_sc_hs__fill_8 FILLER_101_13 ();
 sky130_fd_sc_hs__fill_8 FILLER_101_21 ();
 sky130_fd_sc_hs__fill_8 FILLER_101_29 ();
 sky130_fd_sc_hs__fill_8 FILLER_101_37 ();
 sky130_fd_sc_hs__fill_8 FILLER_101_45 ();
 sky130_fd_sc_hs__fill_4 FILLER_101_53 ();
 sky130_fd_sc_hs__fill_1 FILLER_101_57 ();
 sky130_fd_sc_hs__fill_8 FILLER_101_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_101_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_101_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_101_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_101_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_101_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_101_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_101_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_101_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_101_125 ();
 sky130_fd_sc_hs__fill_2 FILLER_101_133 ();
 sky130_fd_sc_hs__fill_2 FILLER_101_143 ();
 sky130_fd_sc_hs__fill_1 FILLER_101_149 ();
 sky130_fd_sc_hs__fill_4 FILLER_101_156 ();
 sky130_fd_sc_hs__fill_2 FILLER_101_171 ();
 sky130_fd_sc_hs__fill_1 FILLER_101_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_101_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_101_183 ();
 sky130_fd_sc_hs__fill_1 FILLER_101_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_101_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_101_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_101_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_101_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_101_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_101_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_101_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_101_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_101_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_101_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_101_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_101_291 ();
 sky130_fd_sc_hs__fill_4 FILLER_101_299 ();
 sky130_fd_sc_hs__fill_2 FILLER_101_303 ();
 sky130_fd_sc_hs__fill_1 FILLER_101_305 ();
 sky130_fd_sc_hs__fill_8 FILLER_101_340 ();
 sky130_fd_sc_hs__fill_8 FILLER_101_366 ();
 sky130_fd_sc_hs__fill_8 FILLER_101_374 ();
 sky130_fd_sc_hs__fill_8 FILLER_101_382 ();
 sky130_fd_sc_hs__fill_4 FILLER_101_390 ();
 sky130_fd_sc_hs__fill_4 FILLER_101_407 ();
 sky130_fd_sc_hs__fill_2 FILLER_101_411 ();
 sky130_fd_sc_hs__fill_1 FILLER_101_413 ();
 sky130_fd_sc_hs__fill_8 FILLER_101_448 ();
 sky130_fd_sc_hs__fill_2 FILLER_101_456 ();
 sky130_fd_sc_hs__fill_1 FILLER_101_458 ();
 sky130_fd_sc_hs__fill_1 FILLER_101_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_101_492 ();
 sky130_fd_sc_hs__fill_4 FILLER_101_500 ();
 sky130_fd_sc_hs__fill_1 FILLER_101_504 ();
 sky130_fd_sc_hs__fill_4 FILLER_101_508 ();
 sky130_fd_sc_hs__fill_2 FILLER_101_512 ();
 sky130_fd_sc_hs__fill_8 FILLER_101_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_101_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_101_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_102_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_102_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_102_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_102_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_102_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_102_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_102_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_102_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_102_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_102_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_102_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_102_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_102_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_102_88 ();
 sky130_fd_sc_hs__fill_2 FILLER_102_96 ();
 sky130_fd_sc_hs__fill_1 FILLER_102_98 ();
 sky130_fd_sc_hs__fill_2 FILLER_102_131 ();
 sky130_fd_sc_hs__fill_1 FILLER_102_133 ();
 sky130_fd_sc_hs__fill_2 FILLER_102_142 ();
 sky130_fd_sc_hs__fill_1 FILLER_102_144 ();
 sky130_fd_sc_hs__fill_4 FILLER_102_170 ();
 sky130_fd_sc_hs__fill_2 FILLER_102_174 ();
 sky130_fd_sc_hs__fill_1 FILLER_102_176 ();
 sky130_fd_sc_hs__fill_1 FILLER_102_204 ();
 sky130_fd_sc_hs__fill_4 FILLER_102_210 ();
 sky130_fd_sc_hs__fill_1 FILLER_102_214 ();
 sky130_fd_sc_hs__fill_4 FILLER_102_235 ();
 sky130_fd_sc_hs__fill_1 FILLER_102_239 ();
 sky130_fd_sc_hs__fill_8 FILLER_102_269 ();
 sky130_fd_sc_hs__fill_8 FILLER_102_277 ();
 sky130_fd_sc_hs__fill_8 FILLER_102_285 ();
 sky130_fd_sc_hs__fill_8 FILLER_102_293 ();
 sky130_fd_sc_hs__fill_1 FILLER_102_301 ();
 sky130_fd_sc_hs__fill_2 FILLER_102_320 ();
 sky130_fd_sc_hs__fill_1 FILLER_102_322 ();
 sky130_fd_sc_hs__fill_4 FILLER_102_371 ();
 sky130_fd_sc_hs__fill_2 FILLER_102_375 ();
 sky130_fd_sc_hs__fill_8 FILLER_102_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_102_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_102_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_102_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_102_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_102_418 ();
 sky130_fd_sc_hs__fill_4 FILLER_102_426 ();
 sky130_fd_sc_hs__fill_2 FILLER_102_430 ();
 sky130_fd_sc_hs__fill_8 FILLER_102_436 ();
 sky130_fd_sc_hs__fill_1 FILLER_102_444 ();
 sky130_fd_sc_hs__fill_4 FILLER_102_448 ();
 sky130_fd_sc_hs__fill_2 FILLER_102_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_102_477 ();
 sky130_fd_sc_hs__fill_8 FILLER_102_485 ();
 sky130_fd_sc_hs__fill_8 FILLER_102_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_102_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_102_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_102_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_102_526 ();
 sky130_fd_sc_hs__fill_4 FILLER_102_534 ();
 sky130_fd_sc_hs__fill_2 FILLER_102_538 ();
 sky130_fd_sc_hs__fill_4 FILLER_103_0 ();
 sky130_fd_sc_hs__fill_2 FILLER_103_4 ();
 sky130_fd_sc_hs__fill_1 FILLER_103_6 ();
 sky130_fd_sc_hs__fill_8 FILLER_103_15 ();
 sky130_fd_sc_hs__fill_8 FILLER_103_23 ();
 sky130_fd_sc_hs__fill_8 FILLER_103_31 ();
 sky130_fd_sc_hs__fill_8 FILLER_103_39 ();
 sky130_fd_sc_hs__fill_8 FILLER_103_47 ();
 sky130_fd_sc_hs__fill_2 FILLER_103_55 ();
 sky130_fd_sc_hs__fill_1 FILLER_103_57 ();
 sky130_fd_sc_hs__fill_4 FILLER_103_59 ();
 sky130_fd_sc_hs__fill_1 FILLER_103_63 ();
 sky130_fd_sc_hs__fill_8 FILLER_103_73 ();
 sky130_fd_sc_hs__fill_8 FILLER_103_81 ();
 sky130_fd_sc_hs__fill_2 FILLER_103_89 ();
 sky130_fd_sc_hs__fill_8 FILLER_103_108 ();
 sky130_fd_sc_hs__fill_8 FILLER_103_117 ();
 sky130_fd_sc_hs__fill_1 FILLER_103_125 ();
 sky130_fd_sc_hs__fill_2 FILLER_103_129 ();
 sky130_fd_sc_hs__fill_4 FILLER_103_134 ();
 sky130_fd_sc_hs__fill_2 FILLER_103_138 ();
 sky130_fd_sc_hs__fill_2 FILLER_103_155 ();
 sky130_fd_sc_hs__fill_8 FILLER_103_160 ();
 sky130_fd_sc_hs__fill_2 FILLER_103_171 ();
 sky130_fd_sc_hs__fill_1 FILLER_103_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_103_222 ();
 sky130_fd_sc_hs__fill_2 FILLER_103_230 ();
 sky130_fd_sc_hs__fill_2 FILLER_103_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_103_238 ();
 sky130_fd_sc_hs__fill_4 FILLER_103_246 ();
 sky130_fd_sc_hs__fill_4 FILLER_103_255 ();
 sky130_fd_sc_hs__fill_2 FILLER_103_259 ();
 sky130_fd_sc_hs__fill_1 FILLER_103_261 ();
 sky130_fd_sc_hs__fill_2 FILLER_103_265 ();
 sky130_fd_sc_hs__fill_4 FILLER_103_270 ();
 sky130_fd_sc_hs__fill_2 FILLER_103_287 ();
 sky130_fd_sc_hs__fill_1 FILLER_103_289 ();
 sky130_fd_sc_hs__fill_4 FILLER_103_291 ();
 sky130_fd_sc_hs__fill_1 FILLER_103_295 ();
 sky130_fd_sc_hs__fill_8 FILLER_103_334 ();
 sky130_fd_sc_hs__fill_4 FILLER_103_342 ();
 sky130_fd_sc_hs__fill_2 FILLER_103_346 ();
 sky130_fd_sc_hs__fill_8 FILLER_103_349 ();
 sky130_fd_sc_hs__fill_2 FILLER_103_357 ();
 sky130_fd_sc_hs__fill_4 FILLER_103_380 ();
 sky130_fd_sc_hs__fill_1 FILLER_103_384 ();
 sky130_fd_sc_hs__fill_8 FILLER_103_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_103_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_103_423 ();
 sky130_fd_sc_hs__fill_2 FILLER_103_431 ();
 sky130_fd_sc_hs__fill_1 FILLER_103_433 ();
 sky130_fd_sc_hs__fill_8 FILLER_103_443 ();
 sky130_fd_sc_hs__fill_8 FILLER_103_451 ();
 sky130_fd_sc_hs__fill_4 FILLER_103_459 ();
 sky130_fd_sc_hs__fill_1 FILLER_103_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_103_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_103_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_103_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_103_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_103_497 ();
 sky130_fd_sc_hs__fill_1 FILLER_103_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_103_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_103_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_103_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_104_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_104_8 ();
 sky130_fd_sc_hs__fill_4 FILLER_104_16 ();
 sky130_fd_sc_hs__fill_1 FILLER_104_20 ();
 sky130_fd_sc_hs__fill_8 FILLER_104_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_104_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_104_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_104_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_104_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_104_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_104_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_104_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_104_88 ();
 sky130_fd_sc_hs__fill_4 FILLER_104_96 ();
 sky130_fd_sc_hs__fill_2 FILLER_104_140 ();
 sky130_fd_sc_hs__fill_1 FILLER_104_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_104_189 ();
 sky130_fd_sc_hs__fill_4 FILLER_104_197 ();
 sky130_fd_sc_hs__fill_2 FILLER_104_201 ();
 sky130_fd_sc_hs__fill_4 FILLER_104_217 ();
 sky130_fd_sc_hs__fill_4 FILLER_104_244 ();
 sky130_fd_sc_hs__fill_2 FILLER_104_248 ();
 sky130_fd_sc_hs__fill_1 FILLER_104_250 ();
 sky130_fd_sc_hs__fill_4 FILLER_104_275 ();
 sky130_fd_sc_hs__fill_8 FILLER_104_282 ();
 sky130_fd_sc_hs__fill_8 FILLER_104_290 ();
 sky130_fd_sc_hs__fill_8 FILLER_104_298 ();
 sky130_fd_sc_hs__fill_8 FILLER_104_306 ();
 sky130_fd_sc_hs__fill_4 FILLER_104_314 ();
 sky130_fd_sc_hs__fill_1 FILLER_104_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_104_320 ();
 sky130_fd_sc_hs__fill_1 FILLER_104_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_104_350 ();
 sky130_fd_sc_hs__fill_8 FILLER_104_358 ();
 sky130_fd_sc_hs__fill_8 FILLER_104_366 ();
 sky130_fd_sc_hs__fill_2 FILLER_104_374 ();
 sky130_fd_sc_hs__fill_1 FILLER_104_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_104_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_104_386 ();
 sky130_fd_sc_hs__fill_4 FILLER_104_394 ();
 sky130_fd_sc_hs__fill_1 FILLER_104_398 ();
 sky130_fd_sc_hs__fill_8 FILLER_104_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_104_410 ();
 sky130_fd_sc_hs__fill_4 FILLER_104_418 ();
 sky130_fd_sc_hs__fill_2 FILLER_104_422 ();
 sky130_fd_sc_hs__fill_1 FILLER_104_424 ();
 sky130_fd_sc_hs__fill_4 FILLER_104_428 ();
 sky130_fd_sc_hs__fill_2 FILLER_104_432 ();
 sky130_fd_sc_hs__fill_1 FILLER_104_434 ();
 sky130_fd_sc_hs__fill_1 FILLER_104_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_104_443 ();
 sky130_fd_sc_hs__fill_8 FILLER_104_451 ();
 sky130_fd_sc_hs__fill_8 FILLER_104_459 ();
 sky130_fd_sc_hs__fill_8 FILLER_104_467 ();
 sky130_fd_sc_hs__fill_8 FILLER_104_475 ();
 sky130_fd_sc_hs__fill_8 FILLER_104_483 ();
 sky130_fd_sc_hs__fill_2 FILLER_104_491 ();
 sky130_fd_sc_hs__fill_8 FILLER_104_517 ();
 sky130_fd_sc_hs__fill_8 FILLER_104_525 ();
 sky130_fd_sc_hs__fill_4 FILLER_104_533 ();
 sky130_fd_sc_hs__fill_2 FILLER_104_537 ();
 sky130_fd_sc_hs__fill_1 FILLER_104_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_105_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_105_8 ();
 sky130_fd_sc_hs__fill_1 FILLER_105_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_105_25 ();
 sky130_fd_sc_hs__fill_8 FILLER_105_33 ();
 sky130_fd_sc_hs__fill_8 FILLER_105_41 ();
 sky130_fd_sc_hs__fill_8 FILLER_105_49 ();
 sky130_fd_sc_hs__fill_1 FILLER_105_57 ();
 sky130_fd_sc_hs__fill_8 FILLER_105_59 ();
 sky130_fd_sc_hs__fill_1 FILLER_105_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_105_77 ();
 sky130_fd_sc_hs__fill_8 FILLER_105_85 ();
 sky130_fd_sc_hs__fill_8 FILLER_105_93 ();
 sky130_fd_sc_hs__fill_8 FILLER_105_101 ();
 sky130_fd_sc_hs__fill_4 FILLER_105_109 ();
 sky130_fd_sc_hs__fill_2 FILLER_105_113 ();
 sky130_fd_sc_hs__fill_1 FILLER_105_115 ();
 sky130_fd_sc_hs__fill_1 FILLER_105_130 ();
 sky130_fd_sc_hs__fill_8 FILLER_105_155 ();
 sky130_fd_sc_hs__fill_8 FILLER_105_163 ();
 sky130_fd_sc_hs__fill_2 FILLER_105_171 ();
 sky130_fd_sc_hs__fill_1 FILLER_105_173 ();
 sky130_fd_sc_hs__fill_1 FILLER_105_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_105_179 ();
 sky130_fd_sc_hs__fill_8 FILLER_105_187 ();
 sky130_fd_sc_hs__fill_8 FILLER_105_195 ();
 sky130_fd_sc_hs__fill_2 FILLER_105_203 ();
 sky130_fd_sc_hs__fill_8 FILLER_105_210 ();
 sky130_fd_sc_hs__fill_8 FILLER_105_218 ();
 sky130_fd_sc_hs__fill_4 FILLER_105_226 ();
 sky130_fd_sc_hs__fill_2 FILLER_105_230 ();
 sky130_fd_sc_hs__fill_8 FILLER_105_233 ();
 sky130_fd_sc_hs__fill_1 FILLER_105_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_105_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_105_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_105_265 ();
 sky130_fd_sc_hs__fill_1 FILLER_105_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_105_279 ();
 sky130_fd_sc_hs__fill_2 FILLER_105_287 ();
 sky130_fd_sc_hs__fill_1 FILLER_105_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_105_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_105_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_105_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_105_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_105_323 ();
 sky130_fd_sc_hs__fill_4 FILLER_105_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_105_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_105_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_105_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_105_373 ();
 sky130_fd_sc_hs__fill_4 FILLER_105_381 ();
 sky130_fd_sc_hs__fill_2 FILLER_105_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_105_420 ();
 sky130_fd_sc_hs__fill_4 FILLER_105_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_105_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_105_473 ();
 sky130_fd_sc_hs__fill_1 FILLER_105_481 ();
 sky130_fd_sc_hs__fill_4 FILLER_105_518 ();
 sky130_fd_sc_hs__fill_1 FILLER_105_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_106_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_106_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_106_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_106_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_106_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_106_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_106_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_106_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_106_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_106_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_106_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_106_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_106_86 ();
 sky130_fd_sc_hs__fill_4 FILLER_106_88 ();
 sky130_fd_sc_hs__fill_2 FILLER_106_92 ();
 sky130_fd_sc_hs__fill_8 FILLER_106_102 ();
 sky130_fd_sc_hs__fill_8 FILLER_106_110 ();
 sky130_fd_sc_hs__fill_8 FILLER_106_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_106_144 ();
 sky130_fd_sc_hs__fill_4 FILLER_106_146 ();
 sky130_fd_sc_hs__fill_2 FILLER_106_150 ();
 sky130_fd_sc_hs__fill_1 FILLER_106_152 ();
 sky130_fd_sc_hs__fill_8 FILLER_106_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_106_165 ();
 sky130_fd_sc_hs__fill_4 FILLER_106_181 ();
 sky130_fd_sc_hs__fill_1 FILLER_106_185 ();
 sky130_fd_sc_hs__fill_8 FILLER_106_214 ();
 sky130_fd_sc_hs__fill_8 FILLER_106_222 ();
 sky130_fd_sc_hs__fill_8 FILLER_106_230 ();
 sky130_fd_sc_hs__fill_8 FILLER_106_238 ();
 sky130_fd_sc_hs__fill_8 FILLER_106_246 ();
 sky130_fd_sc_hs__fill_4 FILLER_106_254 ();
 sky130_fd_sc_hs__fill_2 FILLER_106_258 ();
 sky130_fd_sc_hs__fill_1 FILLER_106_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_106_262 ();
 sky130_fd_sc_hs__fill_4 FILLER_106_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_106_284 ();
 sky130_fd_sc_hs__fill_4 FILLER_106_292 ();
 sky130_fd_sc_hs__fill_1 FILLER_106_296 ();
 sky130_fd_sc_hs__fill_4 FILLER_106_314 ();
 sky130_fd_sc_hs__fill_1 FILLER_106_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_106_320 ();
 sky130_fd_sc_hs__fill_1 FILLER_106_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_106_345 ();
 sky130_fd_sc_hs__fill_4 FILLER_106_353 ();
 sky130_fd_sc_hs__fill_2 FILLER_106_357 ();
 sky130_fd_sc_hs__fill_1 FILLER_106_359 ();
 sky130_fd_sc_hs__fill_8 FILLER_106_378 ();
 sky130_fd_sc_hs__fill_4 FILLER_106_386 ();
 sky130_fd_sc_hs__fill_2 FILLER_106_390 ();
 sky130_fd_sc_hs__fill_8 FILLER_106_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_106_413 ();
 sky130_fd_sc_hs__fill_4 FILLER_106_421 ();
 sky130_fd_sc_hs__fill_1 FILLER_106_431 ();
 sky130_fd_sc_hs__fill_2 FILLER_106_442 ();
 sky130_fd_sc_hs__fill_8 FILLER_106_467 ();
 sky130_fd_sc_hs__fill_8 FILLER_106_475 ();
 sky130_fd_sc_hs__fill_2 FILLER_106_490 ();
 sky130_fd_sc_hs__fill_1 FILLER_106_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_107_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_107_8 ();
 sky130_fd_sc_hs__fill_1 FILLER_107_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_107_25 ();
 sky130_fd_sc_hs__fill_4 FILLER_107_33 ();
 sky130_fd_sc_hs__fill_2 FILLER_107_37 ();
 sky130_fd_sc_hs__fill_4 FILLER_107_59 ();
 sky130_fd_sc_hs__fill_2 FILLER_107_63 ();
 sky130_fd_sc_hs__fill_1 FILLER_107_65 ();
 sky130_fd_sc_hs__fill_8 FILLER_107_87 ();
 sky130_fd_sc_hs__fill_8 FILLER_107_95 ();
 sky130_fd_sc_hs__fill_8 FILLER_107_103 ();
 sky130_fd_sc_hs__fill_4 FILLER_107_111 ();
 sky130_fd_sc_hs__fill_1 FILLER_107_115 ();
 sky130_fd_sc_hs__fill_4 FILLER_107_129 ();
 sky130_fd_sc_hs__fill_2 FILLER_107_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_107_138 ();
 sky130_fd_sc_hs__fill_8 FILLER_107_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_107_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_107_162 ();
 sky130_fd_sc_hs__fill_4 FILLER_107_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_107_175 ();
 sky130_fd_sc_hs__fill_4 FILLER_107_183 ();
 sky130_fd_sc_hs__fill_4 FILLER_107_190 ();
 sky130_fd_sc_hs__fill_1 FILLER_107_194 ();
 sky130_fd_sc_hs__fill_8 FILLER_107_198 ();
 sky130_fd_sc_hs__fill_8 FILLER_107_206 ();
 sky130_fd_sc_hs__fill_8 FILLER_107_214 ();
 sky130_fd_sc_hs__fill_4 FILLER_107_222 ();
 sky130_fd_sc_hs__fill_2 FILLER_107_229 ();
 sky130_fd_sc_hs__fill_1 FILLER_107_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_107_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_107_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_107_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_107_257 ();
 sky130_fd_sc_hs__fill_4 FILLER_107_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_107_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_107_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_107_307 ();
 sky130_fd_sc_hs__fill_1 FILLER_107_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_107_329 ();
 sky130_fd_sc_hs__fill_8 FILLER_107_337 ();
 sky130_fd_sc_hs__fill_2 FILLER_107_345 ();
 sky130_fd_sc_hs__fill_1 FILLER_107_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_107_349 ();
 sky130_fd_sc_hs__fill_4 FILLER_107_357 ();
 sky130_fd_sc_hs__fill_1 FILLER_107_361 ();
 sky130_fd_sc_hs__fill_8 FILLER_107_375 ();
 sky130_fd_sc_hs__fill_8 FILLER_107_383 ();
 sky130_fd_sc_hs__fill_2 FILLER_107_391 ();
 sky130_fd_sc_hs__fill_1 FILLER_107_393 ();
 sky130_fd_sc_hs__fill_8 FILLER_107_407 ();
 sky130_fd_sc_hs__fill_4 FILLER_107_415 ();
 sky130_fd_sc_hs__fill_4 FILLER_107_443 ();
 sky130_fd_sc_hs__fill_2 FILLER_107_447 ();
 sky130_fd_sc_hs__fill_4 FILLER_107_457 ();
 sky130_fd_sc_hs__fill_2 FILLER_107_461 ();
 sky130_fd_sc_hs__fill_1 FILLER_107_463 ();
 sky130_fd_sc_hs__fill_1 FILLER_107_501 ();
 sky130_fd_sc_hs__fill_1 FILLER_107_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_108_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_108_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_108_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_108_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_108_28 ();
 sky130_fd_sc_hs__fill_2 FILLER_108_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_108_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_108_48 ();
 sky130_fd_sc_hs__fill_8 FILLER_108_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_108_64 ();
 sky130_fd_sc_hs__fill_8 FILLER_108_72 ();
 sky130_fd_sc_hs__fill_4 FILLER_108_80 ();
 sky130_fd_sc_hs__fill_2 FILLER_108_84 ();
 sky130_fd_sc_hs__fill_1 FILLER_108_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_108_113 ();
 sky130_fd_sc_hs__fill_8 FILLER_108_121 ();
 sky130_fd_sc_hs__fill_8 FILLER_108_129 ();
 sky130_fd_sc_hs__fill_2 FILLER_108_137 ();
 sky130_fd_sc_hs__fill_2 FILLER_108_142 ();
 sky130_fd_sc_hs__fill_1 FILLER_108_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_108_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_108_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_108_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_108_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_108_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_108_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_108_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_108_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_108_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_108_212 ();
 sky130_fd_sc_hs__fill_1 FILLER_108_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_108_224 ();
 sky130_fd_sc_hs__fill_1 FILLER_108_232 ();
 sky130_fd_sc_hs__fill_8 FILLER_108_240 ();
 sky130_fd_sc_hs__fill_8 FILLER_108_248 ();
 sky130_fd_sc_hs__fill_4 FILLER_108_256 ();
 sky130_fd_sc_hs__fill_1 FILLER_108_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_108_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_108_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_108_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_108_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_108_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_108_302 ();
 sky130_fd_sc_hs__fill_8 FILLER_108_310 ();
 sky130_fd_sc_hs__fill_1 FILLER_108_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_108_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_108_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_108_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_108_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_108_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_108_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_108_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_108_376 ();
 sky130_fd_sc_hs__fill_2 FILLER_108_378 ();
 sky130_fd_sc_hs__fill_1 FILLER_108_380 ();
 sky130_fd_sc_hs__fill_8 FILLER_108_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_108_413 ();
 sky130_fd_sc_hs__fill_4 FILLER_108_421 ();
 sky130_fd_sc_hs__fill_2 FILLER_108_425 ();
 sky130_fd_sc_hs__fill_1 FILLER_108_427 ();
 sky130_fd_sc_hs__fill_1 FILLER_108_434 ();
 sky130_fd_sc_hs__fill_2 FILLER_108_459 ();
 sky130_fd_sc_hs__fill_8 FILLER_108_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_108_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_108_494 ();
 sky130_fd_sc_hs__fill_1 FILLER_108_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_108_507 ();
 sky130_fd_sc_hs__fill_2 FILLER_108_515 ();
 sky130_fd_sc_hs__fill_1 FILLER_108_517 ();
 sky130_fd_sc_hs__fill_8 FILLER_109_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_109_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_109_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_109_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_109_32 ();
 sky130_fd_sc_hs__fill_2 FILLER_109_41 ();
 sky130_fd_sc_hs__fill_1 FILLER_109_43 ();
 sky130_fd_sc_hs__fill_4 FILLER_109_54 ();
 sky130_fd_sc_hs__fill_2 FILLER_109_59 ();
 sky130_fd_sc_hs__fill_1 FILLER_109_61 ();
 sky130_fd_sc_hs__fill_4 FILLER_109_111 ();
 sky130_fd_sc_hs__fill_1 FILLER_109_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_109_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_109_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_109_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_109_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_109_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_109_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_109_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_109_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_109_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_109_190 ();
 sky130_fd_sc_hs__fill_8 FILLER_109_201 ();
 sky130_fd_sc_hs__fill_1 FILLER_109_209 ();
 sky130_fd_sc_hs__fill_8 FILLER_109_222 ();
 sky130_fd_sc_hs__fill_2 FILLER_109_230 ();
 sky130_fd_sc_hs__fill_8 FILLER_109_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_109_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_109_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_109_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_109_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_109_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_109_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_109_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_109_291 ();
 sky130_fd_sc_hs__fill_2 FILLER_109_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_109_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_109_326 ();
 sky130_fd_sc_hs__fill_8 FILLER_109_334 ();
 sky130_fd_sc_hs__fill_4 FILLER_109_342 ();
 sky130_fd_sc_hs__fill_2 FILLER_109_346 ();
 sky130_fd_sc_hs__fill_4 FILLER_109_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_109_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_109_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_109_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_109_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_109_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_109_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_109_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_109_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_109_423 ();
 sky130_fd_sc_hs__fill_1 FILLER_109_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_109_435 ();
 sky130_fd_sc_hs__fill_8 FILLER_109_443 ();
 sky130_fd_sc_hs__fill_8 FILLER_109_451 ();
 sky130_fd_sc_hs__fill_8 FILLER_109_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_109_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_109_484 ();
 sky130_fd_sc_hs__fill_8 FILLER_109_492 ();
 sky130_fd_sc_hs__fill_4 FILLER_109_500 ();
 sky130_fd_sc_hs__fill_1 FILLER_109_504 ();
 sky130_fd_sc_hs__fill_8 FILLER_109_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_109_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_109_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_109_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_109_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_110_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_110_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_110_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_110_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_110_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_110_30 ();
 sky130_fd_sc_hs__fill_1 FILLER_110_38 ();
 sky130_fd_sc_hs__fill_4 FILLER_110_80 ();
 sky130_fd_sc_hs__fill_2 FILLER_110_84 ();
 sky130_fd_sc_hs__fill_1 FILLER_110_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_110_88 ();
 sky130_fd_sc_hs__fill_2 FILLER_110_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_110_114 ();
 sky130_fd_sc_hs__fill_8 FILLER_110_122 ();
 sky130_fd_sc_hs__fill_8 FILLER_110_130 ();
 sky130_fd_sc_hs__fill_1 FILLER_110_138 ();
 sky130_fd_sc_hs__fill_2 FILLER_110_142 ();
 sky130_fd_sc_hs__fill_1 FILLER_110_144 ();
 sky130_fd_sc_hs__fill_4 FILLER_110_146 ();
 sky130_fd_sc_hs__fill_1 FILLER_110_150 ();
 sky130_fd_sc_hs__fill_8 FILLER_110_159 ();
 sky130_fd_sc_hs__fill_1 FILLER_110_167 ();
 sky130_fd_sc_hs__fill_8 FILLER_110_171 ();
 sky130_fd_sc_hs__fill_1 FILLER_110_182 ();
 sky130_fd_sc_hs__fill_4 FILLER_110_204 ();
 sky130_fd_sc_hs__fill_1 FILLER_110_208 ();
 sky130_fd_sc_hs__fill_4 FILLER_110_219 ();
 sky130_fd_sc_hs__fill_2 FILLER_110_247 ();
 sky130_fd_sc_hs__fill_1 FILLER_110_249 ();
 sky130_fd_sc_hs__fill_2 FILLER_110_253 ();
 sky130_fd_sc_hs__fill_4 FILLER_110_262 ();
 sky130_fd_sc_hs__fill_2 FILLER_110_266 ();
 sky130_fd_sc_hs__fill_1 FILLER_110_268 ();
 sky130_fd_sc_hs__fill_4 FILLER_110_282 ();
 sky130_fd_sc_hs__fill_2 FILLER_110_286 ();
 sky130_fd_sc_hs__fill_2 FILLER_110_295 ();
 sky130_fd_sc_hs__fill_1 FILLER_110_297 ();
 sky130_fd_sc_hs__fill_2 FILLER_110_301 ();
 sky130_fd_sc_hs__fill_4 FILLER_110_320 ();
 sky130_fd_sc_hs__fill_4 FILLER_110_355 ();
 sky130_fd_sc_hs__fill_2 FILLER_110_395 ();
 sky130_fd_sc_hs__fill_8 FILLER_110_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_110_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_110_434 ();
 sky130_fd_sc_hs__fill_2 FILLER_110_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_110_477 ();
 sky130_fd_sc_hs__fill_8 FILLER_110_485 ();
 sky130_fd_sc_hs__fill_8 FILLER_110_494 ();
 sky130_fd_sc_hs__fill_1 FILLER_110_502 ();
 sky130_fd_sc_hs__fill_1 FILLER_110_531 ();
 sky130_fd_sc_hs__fill_2 FILLER_111_0 ();
 sky130_fd_sc_hs__fill_1 FILLER_111_2 ();
 sky130_fd_sc_hs__fill_4 FILLER_111_11 ();
 sky130_fd_sc_hs__fill_1 FILLER_111_15 ();
 sky130_fd_sc_hs__fill_4 FILLER_111_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_111_28 ();
 sky130_fd_sc_hs__fill_4 FILLER_111_41 ();
 sky130_fd_sc_hs__fill_2 FILLER_111_56 ();
 sky130_fd_sc_hs__fill_2 FILLER_111_59 ();
 sky130_fd_sc_hs__fill_1 FILLER_111_61 ();
 sky130_fd_sc_hs__fill_2 FILLER_111_68 ();
 sky130_fd_sc_hs__fill_8 FILLER_111_90 ();
 sky130_fd_sc_hs__fill_8 FILLER_111_98 ();
 sky130_fd_sc_hs__fill_1 FILLER_111_106 ();
 sky130_fd_sc_hs__fill_4 FILLER_111_117 ();
 sky130_fd_sc_hs__fill_1 FILLER_111_121 ();
 sky130_fd_sc_hs__fill_2 FILLER_111_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_111_154 ();
 sky130_fd_sc_hs__fill_4 FILLER_111_162 ();
 sky130_fd_sc_hs__fill_1 FILLER_111_166 ();
 sky130_fd_sc_hs__fill_4 FILLER_111_222 ();
 sky130_fd_sc_hs__fill_2 FILLER_111_226 ();
 sky130_fd_sc_hs__fill_1 FILLER_111_231 ();
 sky130_fd_sc_hs__fill_1 FILLER_111_233 ();
 sky130_fd_sc_hs__fill_1 FILLER_111_237 ();
 sky130_fd_sc_hs__fill_2 FILLER_111_259 ();
 sky130_fd_sc_hs__fill_1 FILLER_111_261 ();
 sky130_fd_sc_hs__fill_8 FILLER_111_268 ();
 sky130_fd_sc_hs__fill_8 FILLER_111_276 ();
 sky130_fd_sc_hs__fill_4 FILLER_111_284 ();
 sky130_fd_sc_hs__fill_2 FILLER_111_288 ();
 sky130_fd_sc_hs__fill_8 FILLER_111_291 ();
 sky130_fd_sc_hs__fill_4 FILLER_111_299 ();
 sky130_fd_sc_hs__fill_1 FILLER_111_303 ();
 sky130_fd_sc_hs__fill_2 FILLER_111_321 ();
 sky130_fd_sc_hs__fill_1 FILLER_111_323 ();
 sky130_fd_sc_hs__fill_4 FILLER_111_328 ();
 sky130_fd_sc_hs__fill_2 FILLER_111_332 ();
 sky130_fd_sc_hs__fill_1 FILLER_111_334 ();
 sky130_fd_sc_hs__fill_8 FILLER_111_349 ();
 sky130_fd_sc_hs__fill_2 FILLER_111_357 ();
 sky130_fd_sc_hs__fill_1 FILLER_111_376 ();
 sky130_fd_sc_hs__fill_1 FILLER_111_380 ();
 sky130_fd_sc_hs__fill_8 FILLER_111_385 ();
 sky130_fd_sc_hs__fill_8 FILLER_111_393 ();
 sky130_fd_sc_hs__fill_4 FILLER_111_401 ();
 sky130_fd_sc_hs__fill_1 FILLER_111_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_111_407 ();
 sky130_fd_sc_hs__fill_1 FILLER_111_415 ();
 sky130_fd_sc_hs__fill_4 FILLER_111_429 ();
 sky130_fd_sc_hs__fill_1 FILLER_111_433 ();
 sky130_fd_sc_hs__fill_4 FILLER_111_454 ();
 sky130_fd_sc_hs__fill_1 FILLER_111_458 ();
 sky130_fd_sc_hs__fill_8 FILLER_111_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_111_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_111_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_111_489 ();
 sky130_fd_sc_hs__fill_4 FILLER_111_497 ();
 sky130_fd_sc_hs__fill_1 FILLER_111_501 ();
 sky130_fd_sc_hs__fill_8 FILLER_111_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_111_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_111_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_112_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_112_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_112_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_112_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_112_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_112_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_112_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_112_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_112_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_112_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_112_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_112_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_112_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_112_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_112_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_112_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_112_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_112_120 ();
 sky130_fd_sc_hs__fill_2 FILLER_112_128 ();
 sky130_fd_sc_hs__fill_2 FILLER_112_143 ();
 sky130_fd_sc_hs__fill_8 FILLER_112_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_112_154 ();
 sky130_fd_sc_hs__fill_4 FILLER_112_162 ();
 sky130_fd_sc_hs__fill_2 FILLER_112_166 ();
 sky130_fd_sc_hs__fill_1 FILLER_112_172 ();
 sky130_fd_sc_hs__fill_8 FILLER_112_180 ();
 sky130_fd_sc_hs__fill_2 FILLER_112_188 ();
 sky130_fd_sc_hs__fill_8 FILLER_112_193 ();
 sky130_fd_sc_hs__fill_2 FILLER_112_201 ();
 sky130_fd_sc_hs__fill_1 FILLER_112_204 ();
 sky130_fd_sc_hs__fill_4 FILLER_112_239 ();
 sky130_fd_sc_hs__fill_1 FILLER_112_243 ();
 sky130_fd_sc_hs__fill_2 FILLER_112_247 ();
 sky130_fd_sc_hs__fill_2 FILLER_112_256 ();
 sky130_fd_sc_hs__fill_8 FILLER_112_283 ();
 sky130_fd_sc_hs__fill_8 FILLER_112_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_112_299 ();
 sky130_fd_sc_hs__fill_2 FILLER_112_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_112_320 ();
 sky130_fd_sc_hs__fill_4 FILLER_112_344 ();
 sky130_fd_sc_hs__fill_2 FILLER_112_348 ();
 sky130_fd_sc_hs__fill_1 FILLER_112_350 ();
 sky130_fd_sc_hs__fill_4 FILLER_112_372 ();
 sky130_fd_sc_hs__fill_1 FILLER_112_376 ();
 sky130_fd_sc_hs__fill_4 FILLER_112_398 ();
 sky130_fd_sc_hs__fill_2 FILLER_112_402 ();
 sky130_fd_sc_hs__fill_1 FILLER_112_404 ();
 sky130_fd_sc_hs__fill_4 FILLER_112_436 ();
 sky130_fd_sc_hs__fill_2 FILLER_112_440 ();
 sky130_fd_sc_hs__fill_1 FILLER_112_442 ();
 sky130_fd_sc_hs__fill_2 FILLER_112_487 ();
 sky130_fd_sc_hs__fill_1 FILLER_112_489 ();
 sky130_fd_sc_hs__fill_1 FILLER_112_494 ();
 sky130_fd_sc_hs__fill_1 FILLER_112_499 ();
 sky130_fd_sc_hs__fill_2 FILLER_112_538 ();
 sky130_fd_sc_hs__fill_8 FILLER_113_0 ();
 sky130_fd_sc_hs__fill_4 FILLER_113_8 ();
 sky130_fd_sc_hs__fill_1 FILLER_113_12 ();
 sky130_fd_sc_hs__fill_8 FILLER_113_21 ();
 sky130_fd_sc_hs__fill_8 FILLER_113_29 ();
 sky130_fd_sc_hs__fill_2 FILLER_113_37 ();
 sky130_fd_sc_hs__fill_4 FILLER_113_52 ();
 sky130_fd_sc_hs__fill_2 FILLER_113_56 ();
 sky130_fd_sc_hs__fill_2 FILLER_113_59 ();
 sky130_fd_sc_hs__fill_1 FILLER_113_61 ();
 sky130_fd_sc_hs__fill_8 FILLER_113_93 ();
 sky130_fd_sc_hs__fill_8 FILLER_113_101 ();
 sky130_fd_sc_hs__fill_4 FILLER_113_109 ();
 sky130_fd_sc_hs__fill_2 FILLER_113_113 ();
 sky130_fd_sc_hs__fill_1 FILLER_113_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_113_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_113_152 ();
 sky130_fd_sc_hs__fill_8 FILLER_113_160 ();
 sky130_fd_sc_hs__fill_4 FILLER_113_168 ();
 sky130_fd_sc_hs__fill_2 FILLER_113_172 ();
 sky130_fd_sc_hs__fill_4 FILLER_113_175 ();
 sky130_fd_sc_hs__fill_2 FILLER_113_179 ();
 sky130_fd_sc_hs__fill_1 FILLER_113_181 ();
 sky130_fd_sc_hs__fill_8 FILLER_113_189 ();
 sky130_fd_sc_hs__fill_2 FILLER_113_197 ();
 sky130_fd_sc_hs__fill_4 FILLER_113_202 ();
 sky130_fd_sc_hs__fill_2 FILLER_113_206 ();
 sky130_fd_sc_hs__fill_1 FILLER_113_214 ();
 sky130_fd_sc_hs__fill_8 FILLER_113_222 ();
 sky130_fd_sc_hs__fill_2 FILLER_113_230 ();
 sky130_fd_sc_hs__fill_8 FILLER_113_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_113_241 ();
 sky130_fd_sc_hs__fill_2 FILLER_113_249 ();
 sky130_fd_sc_hs__fill_1 FILLER_113_251 ();
 sky130_fd_sc_hs__fill_8 FILLER_113_255 ();
 sky130_fd_sc_hs__fill_2 FILLER_113_270 ();
 sky130_fd_sc_hs__fill_1 FILLER_113_272 ();
 sky130_fd_sc_hs__fill_8 FILLER_113_280 ();
 sky130_fd_sc_hs__fill_2 FILLER_113_288 ();
 sky130_fd_sc_hs__fill_8 FILLER_113_291 ();
 sky130_fd_sc_hs__fill_4 FILLER_113_299 ();
 sky130_fd_sc_hs__fill_2 FILLER_113_303 ();
 sky130_fd_sc_hs__fill_1 FILLER_113_305 ();
 sky130_fd_sc_hs__fill_8 FILLER_113_316 ();
 sky130_fd_sc_hs__fill_4 FILLER_113_324 ();
 sky130_fd_sc_hs__fill_8 FILLER_113_338 ();
 sky130_fd_sc_hs__fill_2 FILLER_113_346 ();
 sky130_fd_sc_hs__fill_8 FILLER_113_349 ();
 sky130_fd_sc_hs__fill_4 FILLER_113_357 ();
 sky130_fd_sc_hs__fill_1 FILLER_113_361 ();
 sky130_fd_sc_hs__fill_8 FILLER_113_375 ();
 sky130_fd_sc_hs__fill_8 FILLER_113_383 ();
 sky130_fd_sc_hs__fill_8 FILLER_113_391 ();
 sky130_fd_sc_hs__fill_4 FILLER_113_399 ();
 sky130_fd_sc_hs__fill_2 FILLER_113_403 ();
 sky130_fd_sc_hs__fill_1 FILLER_113_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_113_424 ();
 sky130_fd_sc_hs__fill_8 FILLER_113_432 ();
 sky130_fd_sc_hs__fill_8 FILLER_113_440 ();
 sky130_fd_sc_hs__fill_8 FILLER_113_448 ();
 sky130_fd_sc_hs__fill_8 FILLER_113_456 ();
 sky130_fd_sc_hs__fill_8 FILLER_113_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_113_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_113_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_113_489 ();
 sky130_fd_sc_hs__fill_2 FILLER_113_520 ();
 sky130_fd_sc_hs__fill_2 FILLER_113_529 ();
 sky130_fd_sc_hs__fill_1 FILLER_113_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_114_0 ();
 sky130_fd_sc_hs__fill_4 FILLER_114_8 ();
 sky130_fd_sc_hs__fill_1 FILLER_114_12 ();
 sky130_fd_sc_hs__fill_8 FILLER_114_21 ();
 sky130_fd_sc_hs__fill_8 FILLER_114_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_114_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_114_46 ();
 sky130_fd_sc_hs__fill_4 FILLER_114_54 ();
 sky130_fd_sc_hs__fill_1 FILLER_114_58 ();
 sky130_fd_sc_hs__fill_8 FILLER_114_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_114_96 ();
 sky130_fd_sc_hs__fill_4 FILLER_114_104 ();
 sky130_fd_sc_hs__fill_2 FILLER_114_108 ();
 sky130_fd_sc_hs__fill_4 FILLER_114_124 ();
 sky130_fd_sc_hs__fill_8 FILLER_114_154 ();
 sky130_fd_sc_hs__fill_2 FILLER_114_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_114_179 ();
 sky130_fd_sc_hs__fill_8 FILLER_114_187 ();
 sky130_fd_sc_hs__fill_4 FILLER_114_195 ();
 sky130_fd_sc_hs__fill_8 FILLER_114_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_114_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_114_220 ();
 sky130_fd_sc_hs__fill_1 FILLER_114_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_114_237 ();
 sky130_fd_sc_hs__fill_8 FILLER_114_245 ();
 sky130_fd_sc_hs__fill_8 FILLER_114_253 ();
 sky130_fd_sc_hs__fill_8 FILLER_114_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_114_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_114_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_114_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_114_294 ();
 sky130_fd_sc_hs__fill_2 FILLER_114_302 ();
 sky130_fd_sc_hs__fill_1 FILLER_114_304 ();
 sky130_fd_sc_hs__fill_8 FILLER_114_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_114_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_114_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_114_361 ();
 sky130_fd_sc_hs__fill_8 FILLER_114_369 ();
 sky130_fd_sc_hs__fill_8 FILLER_114_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_114_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_114_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_114_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_114_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_114_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_114_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_114_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_114_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_114_444 ();
 sky130_fd_sc_hs__fill_4 FILLER_114_452 ();
 sky130_fd_sc_hs__fill_2 FILLER_114_456 ();
 sky130_fd_sc_hs__fill_8 FILLER_114_482 ();
 sky130_fd_sc_hs__fill_2 FILLER_114_490 ();
 sky130_fd_sc_hs__fill_1 FILLER_114_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_114_494 ();
 sky130_fd_sc_hs__fill_4 FILLER_114_502 ();
 sky130_fd_sc_hs__fill_2 FILLER_114_506 ();
 sky130_fd_sc_hs__fill_1 FILLER_114_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_115_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_115_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_115_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_115_24 ();
 sky130_fd_sc_hs__fill_4 FILLER_115_32 ();
 sky130_fd_sc_hs__fill_1 FILLER_115_57 ();
 sky130_fd_sc_hs__fill_4 FILLER_115_59 ();
 sky130_fd_sc_hs__fill_1 FILLER_115_63 ();
 sky130_fd_sc_hs__fill_8 FILLER_115_82 ();
 sky130_fd_sc_hs__fill_8 FILLER_115_90 ();
 sky130_fd_sc_hs__fill_8 FILLER_115_98 ();
 sky130_fd_sc_hs__fill_8 FILLER_115_106 ();
 sky130_fd_sc_hs__fill_2 FILLER_115_114 ();
 sky130_fd_sc_hs__fill_8 FILLER_115_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_115_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_115_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_115_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_115_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_115_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_115_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_115_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_115_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_115_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_115_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_115_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_115_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_115_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_115_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_115_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_115_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_115_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_115_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_115_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_115_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_115_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_115_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_115_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_115_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_115_299 ();
 sky130_fd_sc_hs__fill_4 FILLER_115_307 ();
 sky130_fd_sc_hs__fill_2 FILLER_115_311 ();
 sky130_fd_sc_hs__fill_1 FILLER_115_313 ();
 sky130_fd_sc_hs__fill_8 FILLER_115_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_115_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_115_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_115_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_115_357 ();
 sky130_fd_sc_hs__fill_2 FILLER_115_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_115_375 ();
 sky130_fd_sc_hs__fill_8 FILLER_115_383 ();
 sky130_fd_sc_hs__fill_4 FILLER_115_391 ();
 sky130_fd_sc_hs__fill_2 FILLER_115_395 ();
 sky130_fd_sc_hs__fill_8 FILLER_115_407 ();
 sky130_fd_sc_hs__fill_2 FILLER_115_415 ();
 sky130_fd_sc_hs__fill_1 FILLER_115_417 ();
 sky130_fd_sc_hs__fill_8 FILLER_115_435 ();
 sky130_fd_sc_hs__fill_8 FILLER_115_443 ();
 sky130_fd_sc_hs__fill_4 FILLER_115_451 ();
 sky130_fd_sc_hs__fill_1 FILLER_115_455 ();
 sky130_fd_sc_hs__fill_4 FILLER_115_459 ();
 sky130_fd_sc_hs__fill_1 FILLER_115_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_115_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_115_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_115_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_115_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_115_497 ();
 sky130_fd_sc_hs__fill_1 FILLER_115_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_115_514 ();
 sky130_fd_sc_hs__fill_8 FILLER_115_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_115_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_115_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_116_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_116_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_116_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_116_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_116_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_116_30 ();
 sky130_fd_sc_hs__fill_4 FILLER_116_38 ();
 sky130_fd_sc_hs__fill_1 FILLER_116_42 ();
 sky130_fd_sc_hs__fill_8 FILLER_116_61 ();
 sky130_fd_sc_hs__fill_8 FILLER_116_69 ();
 sky130_fd_sc_hs__fill_8 FILLER_116_77 ();
 sky130_fd_sc_hs__fill_2 FILLER_116_85 ();
 sky130_fd_sc_hs__fill_8 FILLER_116_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_116_96 ();
 sky130_fd_sc_hs__fill_2 FILLER_116_104 ();
 sky130_fd_sc_hs__fill_4 FILLER_116_115 ();
 sky130_fd_sc_hs__fill_2 FILLER_116_119 ();
 sky130_fd_sc_hs__fill_1 FILLER_116_121 ();
 sky130_fd_sc_hs__fill_8 FILLER_116_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_116_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_116_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_116_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_116_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_116_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_116_178 ();
 sky130_fd_sc_hs__fill_2 FILLER_116_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_116_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_116_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_116_223 ();
 sky130_fd_sc_hs__fill_8 FILLER_116_231 ();
 sky130_fd_sc_hs__fill_1 FILLER_116_239 ();
 sky130_fd_sc_hs__fill_4 FILLER_116_254 ();
 sky130_fd_sc_hs__fill_8 FILLER_116_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_116_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_116_281 ();
 sky130_fd_sc_hs__fill_8 FILLER_116_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_116_310 ();
 sky130_fd_sc_hs__fill_1 FILLER_116_318 ();
 sky130_fd_sc_hs__fill_4 FILLER_116_320 ();
 sky130_fd_sc_hs__fill_2 FILLER_116_324 ();
 sky130_fd_sc_hs__fill_8 FILLER_116_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_116_352 ();
 sky130_fd_sc_hs__fill_4 FILLER_116_360 ();
 sky130_fd_sc_hs__fill_1 FILLER_116_364 ();
 sky130_fd_sc_hs__fill_8 FILLER_116_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_116_386 ();
 sky130_fd_sc_hs__fill_2 FILLER_116_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_116_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_116_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_116_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_116_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_116_444 ();
 sky130_fd_sc_hs__fill_4 FILLER_116_452 ();
 sky130_fd_sc_hs__fill_1 FILLER_116_456 ();
 sky130_fd_sc_hs__fill_1 FILLER_116_464 ();
 sky130_fd_sc_hs__fill_8 FILLER_116_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_116_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_116_510 ();
 sky130_fd_sc_hs__fill_1 FILLER_116_518 ();
 sky130_fd_sc_hs__fill_4 FILLER_117_0 ();
 sky130_fd_sc_hs__fill_1 FILLER_117_4 ();
 sky130_fd_sc_hs__fill_8 FILLER_117_13 ();
 sky130_fd_sc_hs__fill_8 FILLER_117_29 ();
 sky130_fd_sc_hs__fill_8 FILLER_117_37 ();
 sky130_fd_sc_hs__fill_8 FILLER_117_45 ();
 sky130_fd_sc_hs__fill_4 FILLER_117_53 ();
 sky130_fd_sc_hs__fill_1 FILLER_117_57 ();
 sky130_fd_sc_hs__fill_8 FILLER_117_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_117_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_117_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_117_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_117_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_117_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_117_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_117_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_117_141 ();
 sky130_fd_sc_hs__fill_4 FILLER_117_149 ();
 sky130_fd_sc_hs__fill_2 FILLER_117_153 ();
 sky130_fd_sc_hs__fill_8 FILLER_117_158 ();
 sky130_fd_sc_hs__fill_2 FILLER_117_166 ();
 sky130_fd_sc_hs__fill_2 FILLER_117_171 ();
 sky130_fd_sc_hs__fill_1 FILLER_117_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_117_175 ();
 sky130_fd_sc_hs__fill_4 FILLER_117_183 ();
 sky130_fd_sc_hs__fill_1 FILLER_117_187 ();
 sky130_fd_sc_hs__fill_1 FILLER_117_218 ();
 sky130_fd_sc_hs__fill_2 FILLER_117_226 ();
 sky130_fd_sc_hs__fill_2 FILLER_117_243 ();
 sky130_fd_sc_hs__fill_1 FILLER_117_249 ();
 sky130_fd_sc_hs__fill_4 FILLER_117_258 ();
 sky130_fd_sc_hs__fill_2 FILLER_117_262 ();
 sky130_fd_sc_hs__fill_1 FILLER_117_264 ();
 sky130_fd_sc_hs__fill_8 FILLER_117_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_117_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_117_289 ();
 sky130_fd_sc_hs__fill_2 FILLER_117_291 ();
 sky130_fd_sc_hs__fill_4 FILLER_117_306 ();
 sky130_fd_sc_hs__fill_4 FILLER_117_316 ();
 sky130_fd_sc_hs__fill_2 FILLER_117_320 ();
 sky130_fd_sc_hs__fill_4 FILLER_117_332 ();
 sky130_fd_sc_hs__fill_2 FILLER_117_336 ();
 sky130_fd_sc_hs__fill_1 FILLER_117_359 ();
 sky130_fd_sc_hs__fill_8 FILLER_117_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_117_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_117_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_117_407 ();
 sky130_fd_sc_hs__fill_2 FILLER_117_415 ();
 sky130_fd_sc_hs__fill_1 FILLER_117_450 ();
 sky130_fd_sc_hs__fill_4 FILLER_117_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_117_485 ();
 sky130_fd_sc_hs__fill_8 FILLER_117_493 ();
 sky130_fd_sc_hs__fill_8 FILLER_117_501 ();
 sky130_fd_sc_hs__fill_8 FILLER_117_509 ();
 sky130_fd_sc_hs__fill_4 FILLER_117_517 ();
 sky130_fd_sc_hs__fill_1 FILLER_117_521 ();
 sky130_fd_sc_hs__fill_4 FILLER_117_523 ();
 sky130_fd_sc_hs__fill_4 FILLER_117_535 ();
 sky130_fd_sc_hs__fill_1 FILLER_117_539 ();
 sky130_fd_sc_hs__fill_1 FILLER_118_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_118_9 ();
 sky130_fd_sc_hs__fill_8 FILLER_118_17 ();
 sky130_fd_sc_hs__fill_4 FILLER_118_25 ();
 sky130_fd_sc_hs__fill_8 FILLER_118_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_118_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_118_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_118_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_118_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_118_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_118_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_118_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_118_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_118_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_118_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_118_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_118_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_118_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_118_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_118_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_118_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_118_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_118_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_118_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_118_178 ();
 sky130_fd_sc_hs__fill_1 FILLER_118_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_118_191 ();
 sky130_fd_sc_hs__fill_4 FILLER_118_199 ();
 sky130_fd_sc_hs__fill_2 FILLER_118_204 ();
 sky130_fd_sc_hs__fill_4 FILLER_118_234 ();
 sky130_fd_sc_hs__fill_2 FILLER_118_238 ();
 sky130_fd_sc_hs__fill_8 FILLER_118_243 ();
 sky130_fd_sc_hs__fill_8 FILLER_118_251 ();
 sky130_fd_sc_hs__fill_2 FILLER_118_259 ();
 sky130_fd_sc_hs__fill_4 FILLER_118_262 ();
 sky130_fd_sc_hs__fill_1 FILLER_118_266 ();
 sky130_fd_sc_hs__fill_8 FILLER_118_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_118_281 ();
 sky130_fd_sc_hs__fill_8 FILLER_118_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_118_297 ();
 sky130_fd_sc_hs__fill_4 FILLER_118_305 ();
 sky130_fd_sc_hs__fill_2 FILLER_118_309 ();
 sky130_fd_sc_hs__fill_1 FILLER_118_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_118_339 ();
 sky130_fd_sc_hs__fill_8 FILLER_118_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_118_355 ();
 sky130_fd_sc_hs__fill_4 FILLER_118_363 ();
 sky130_fd_sc_hs__fill_1 FILLER_118_367 ();
 sky130_fd_sc_hs__fill_1 FILLER_118_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_118_378 ();
 sky130_fd_sc_hs__fill_4 FILLER_118_386 ();
 sky130_fd_sc_hs__fill_1 FILLER_118_390 ();
 sky130_fd_sc_hs__fill_8 FILLER_118_413 ();
 sky130_fd_sc_hs__fill_8 FILLER_118_421 ();
 sky130_fd_sc_hs__fill_4 FILLER_118_429 ();
 sky130_fd_sc_hs__fill_2 FILLER_118_433 ();
 sky130_fd_sc_hs__fill_1 FILLER_118_436 ();
 sky130_fd_sc_hs__fill_2 FILLER_118_473 ();
 sky130_fd_sc_hs__fill_1 FILLER_118_475 ();
 sky130_fd_sc_hs__fill_8 FILLER_118_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_118_502 ();
 sky130_fd_sc_hs__fill_2 FILLER_118_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_118_532 ();
 sky130_fd_sc_hs__fill_8 FILLER_119_0 ();
 sky130_fd_sc_hs__fill_4 FILLER_119_8 ();
 sky130_fd_sc_hs__fill_1 FILLER_119_12 ();
 sky130_fd_sc_hs__fill_8 FILLER_119_21 ();
 sky130_fd_sc_hs__fill_8 FILLER_119_29 ();
 sky130_fd_sc_hs__fill_8 FILLER_119_37 ();
 sky130_fd_sc_hs__fill_8 FILLER_119_45 ();
 sky130_fd_sc_hs__fill_4 FILLER_119_53 ();
 sky130_fd_sc_hs__fill_1 FILLER_119_57 ();
 sky130_fd_sc_hs__fill_4 FILLER_119_59 ();
 sky130_fd_sc_hs__fill_2 FILLER_119_63 ();
 sky130_fd_sc_hs__fill_1 FILLER_119_65 ();
 sky130_fd_sc_hs__fill_4 FILLER_119_71 ();
 sky130_fd_sc_hs__fill_8 FILLER_119_78 ();
 sky130_fd_sc_hs__fill_8 FILLER_119_86 ();
 sky130_fd_sc_hs__fill_4 FILLER_119_94 ();
 sky130_fd_sc_hs__fill_2 FILLER_119_98 ();
 sky130_fd_sc_hs__fill_1 FILLER_119_100 ();
 sky130_fd_sc_hs__fill_8 FILLER_119_108 ();
 sky130_fd_sc_hs__fill_8 FILLER_119_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_119_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_119_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_119_141 ();
 sky130_fd_sc_hs__fill_4 FILLER_119_149 ();
 sky130_fd_sc_hs__fill_2 FILLER_119_153 ();
 sky130_fd_sc_hs__fill_1 FILLER_119_155 ();
 sky130_fd_sc_hs__fill_4 FILLER_119_164 ();
 sky130_fd_sc_hs__fill_1 FILLER_119_168 ();
 sky130_fd_sc_hs__fill_4 FILLER_119_184 ();
 sky130_fd_sc_hs__fill_2 FILLER_119_188 ();
 sky130_fd_sc_hs__fill_1 FILLER_119_190 ();
 sky130_fd_sc_hs__fill_2 FILLER_119_198 ();
 sky130_fd_sc_hs__fill_1 FILLER_119_200 ();
 sky130_fd_sc_hs__fill_8 FILLER_119_206 ();
 sky130_fd_sc_hs__fill_8 FILLER_119_214 ();
 sky130_fd_sc_hs__fill_1 FILLER_119_222 ();
 sky130_fd_sc_hs__fill_2 FILLER_119_226 ();
 sky130_fd_sc_hs__fill_1 FILLER_119_228 ();
 sky130_fd_sc_hs__fill_4 FILLER_119_254 ();
 sky130_fd_sc_hs__fill_2 FILLER_119_258 ();
 sky130_fd_sc_hs__fill_1 FILLER_119_260 ();
 sky130_fd_sc_hs__fill_1 FILLER_119_264 ();
 sky130_fd_sc_hs__fill_8 FILLER_119_271 ();
 sky130_fd_sc_hs__fill_8 FILLER_119_279 ();
 sky130_fd_sc_hs__fill_2 FILLER_119_287 ();
 sky130_fd_sc_hs__fill_1 FILLER_119_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_119_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_119_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_119_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_119_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_119_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_119_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_119_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_119_347 ();
 sky130_fd_sc_hs__fill_2 FILLER_119_349 ();
 sky130_fd_sc_hs__fill_1 FILLER_119_351 ();
 sky130_fd_sc_hs__fill_8 FILLER_119_361 ();
 sky130_fd_sc_hs__fill_2 FILLER_119_378 ();
 sky130_fd_sc_hs__fill_1 FILLER_119_380 ();
 sky130_fd_sc_hs__fill_4 FILLER_119_386 ();
 sky130_fd_sc_hs__fill_2 FILLER_119_395 ();
 sky130_fd_sc_hs__fill_8 FILLER_119_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_119_415 ();
 sky130_fd_sc_hs__fill_4 FILLER_119_423 ();
 sky130_fd_sc_hs__fill_2 FILLER_119_427 ();
 sky130_fd_sc_hs__fill_8 FILLER_119_436 ();
 sky130_fd_sc_hs__fill_4 FILLER_119_444 ();
 sky130_fd_sc_hs__fill_1 FILLER_119_448 ();
 sky130_fd_sc_hs__fill_2 FILLER_119_462 ();
 sky130_fd_sc_hs__fill_4 FILLER_119_465 ();
 sky130_fd_sc_hs__fill_2 FILLER_119_469 ();
 sky130_fd_sc_hs__fill_2 FILLER_119_474 ();
 sky130_fd_sc_hs__fill_1 FILLER_119_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_119_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_119_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_119_505 ();
 sky130_fd_sc_hs__fill_2 FILLER_119_519 ();
 sky130_fd_sc_hs__fill_1 FILLER_119_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_119_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_119_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_119_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_120_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_120_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_120_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_120_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_120_28 ();
 sky130_fd_sc_hs__fill_4 FILLER_120_30 ();
 sky130_fd_sc_hs__fill_2 FILLER_120_34 ();
 sky130_fd_sc_hs__fill_2 FILLER_120_41 ();
 sky130_fd_sc_hs__fill_1 FILLER_120_43 ();
 sky130_fd_sc_hs__fill_1 FILLER_120_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_120_88 ();
 sky130_fd_sc_hs__fill_4 FILLER_120_96 ();
 sky130_fd_sc_hs__fill_1 FILLER_120_100 ();
 sky130_fd_sc_hs__fill_8 FILLER_120_146 ();
 sky130_fd_sc_hs__fill_4 FILLER_120_154 ();
 sky130_fd_sc_hs__fill_1 FILLER_120_158 ();
 sky130_fd_sc_hs__fill_8 FILLER_120_180 ();
 sky130_fd_sc_hs__fill_1 FILLER_120_188 ();
 sky130_fd_sc_hs__fill_1 FILLER_120_192 ();
 sky130_fd_sc_hs__fill_1 FILLER_120_196 ();
 sky130_fd_sc_hs__fill_4 FILLER_120_204 ();
 sky130_fd_sc_hs__fill_1 FILLER_120_208 ();
 sky130_fd_sc_hs__fill_8 FILLER_120_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_120_220 ();
 sky130_fd_sc_hs__fill_4 FILLER_120_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_120_243 ();
 sky130_fd_sc_hs__fill_4 FILLER_120_251 ();
 sky130_fd_sc_hs__fill_1 FILLER_120_255 ();
 sky130_fd_sc_hs__fill_2 FILLER_120_259 ();
 sky130_fd_sc_hs__fill_1 FILLER_120_283 ();
 sky130_fd_sc_hs__fill_8 FILLER_120_301 ();
 sky130_fd_sc_hs__fill_8 FILLER_120_309 ();
 sky130_fd_sc_hs__fill_2 FILLER_120_317 ();
 sky130_fd_sc_hs__fill_8 FILLER_120_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_120_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_120_336 ();
 sky130_fd_sc_hs__fill_4 FILLER_120_344 ();
 sky130_fd_sc_hs__fill_2 FILLER_120_348 ();
 sky130_fd_sc_hs__fill_1 FILLER_120_350 ();
 sky130_fd_sc_hs__fill_4 FILLER_120_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_120_400 ();
 sky130_fd_sc_hs__fill_8 FILLER_120_408 ();
 sky130_fd_sc_hs__fill_2 FILLER_120_416 ();
 sky130_fd_sc_hs__fill_8 FILLER_120_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_120_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_120_452 ();
 sky130_fd_sc_hs__fill_1 FILLER_120_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_120_469 ();
 sky130_fd_sc_hs__fill_4 FILLER_120_477 ();
 sky130_fd_sc_hs__fill_8 FILLER_120_494 ();
 sky130_fd_sc_hs__fill_4 FILLER_120_502 ();
 sky130_fd_sc_hs__fill_2 FILLER_120_506 ();
 sky130_fd_sc_hs__fill_1 FILLER_120_516 ();
 sky130_fd_sc_hs__fill_8 FILLER_120_525 ();
 sky130_fd_sc_hs__fill_4 FILLER_120_533 ();
 sky130_fd_sc_hs__fill_2 FILLER_120_537 ();
 sky130_fd_sc_hs__fill_1 FILLER_120_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_121_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_121_8 ();
 sky130_fd_sc_hs__fill_1 FILLER_121_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_121_25 ();
 sky130_fd_sc_hs__fill_8 FILLER_121_45 ();
 sky130_fd_sc_hs__fill_4 FILLER_121_53 ();
 sky130_fd_sc_hs__fill_1 FILLER_121_57 ();
 sky130_fd_sc_hs__fill_2 FILLER_121_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_121_94 ();
 sky130_fd_sc_hs__fill_8 FILLER_121_102 ();
 sky130_fd_sc_hs__fill_4 FILLER_121_110 ();
 sky130_fd_sc_hs__fill_2 FILLER_121_114 ();
 sky130_fd_sc_hs__fill_8 FILLER_121_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_121_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_121_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_121_141 ();
 sky130_fd_sc_hs__fill_2 FILLER_121_149 ();
 sky130_fd_sc_hs__fill_1 FILLER_121_151 ();
 sky130_fd_sc_hs__fill_4 FILLER_121_168 ();
 sky130_fd_sc_hs__fill_2 FILLER_121_172 ();
 sky130_fd_sc_hs__fill_8 FILLER_121_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_121_183 ();
 sky130_fd_sc_hs__fill_4 FILLER_121_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_121_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_121_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_121_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_121_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_121_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_121_244 ();
 sky130_fd_sc_hs__fill_4 FILLER_121_252 ();
 sky130_fd_sc_hs__fill_4 FILLER_121_277 ();
 sky130_fd_sc_hs__fill_8 FILLER_121_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_121_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_121_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_121_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_121_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_121_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_121_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_121_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_121_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_121_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_121_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_121_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_121_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_121_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_121_415 ();
 sky130_fd_sc_hs__fill_1 FILLER_121_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_121_427 ();
 sky130_fd_sc_hs__fill_8 FILLER_121_435 ();
 sky130_fd_sc_hs__fill_8 FILLER_121_443 ();
 sky130_fd_sc_hs__fill_8 FILLER_121_451 ();
 sky130_fd_sc_hs__fill_4 FILLER_121_459 ();
 sky130_fd_sc_hs__fill_1 FILLER_121_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_121_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_121_473 ();
 sky130_fd_sc_hs__fill_4 FILLER_121_481 ();
 sky130_fd_sc_hs__fill_1 FILLER_121_485 ();
 sky130_fd_sc_hs__fill_8 FILLER_121_504 ();
 sky130_fd_sc_hs__fill_8 FILLER_121_512 ();
 sky130_fd_sc_hs__fill_2 FILLER_121_520 ();
 sky130_fd_sc_hs__fill_1 FILLER_121_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_121_532 ();
 sky130_fd_sc_hs__fill_4 FILLER_122_0 ();
 sky130_fd_sc_hs__fill_1 FILLER_122_4 ();
 sky130_fd_sc_hs__fill_8 FILLER_122_13 ();
 sky130_fd_sc_hs__fill_8 FILLER_122_21 ();
 sky130_fd_sc_hs__fill_2 FILLER_122_30 ();
 sky130_fd_sc_hs__fill_1 FILLER_122_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_122_51 ();
 sky130_fd_sc_hs__fill_4 FILLER_122_59 ();
 sky130_fd_sc_hs__fill_2 FILLER_122_63 ();
 sky130_fd_sc_hs__fill_4 FILLER_122_74 ();
 sky130_fd_sc_hs__fill_4 FILLER_122_83 ();
 sky130_fd_sc_hs__fill_4 FILLER_122_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_122_126 ();
 sky130_fd_sc_hs__fill_2 FILLER_122_134 ();
 sky130_fd_sc_hs__fill_1 FILLER_122_136 ();
 sky130_fd_sc_hs__fill_4 FILLER_122_140 ();
 sky130_fd_sc_hs__fill_1 FILLER_122_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_122_146 ();
 sky130_fd_sc_hs__fill_2 FILLER_122_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_122_169 ();
 sky130_fd_sc_hs__fill_4 FILLER_122_177 ();
 sky130_fd_sc_hs__fill_1 FILLER_122_181 ();
 sky130_fd_sc_hs__fill_8 FILLER_122_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_122_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_122_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_122_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_122_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_122_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_122_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_122_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_122_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_122_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_122_278 ();
 sky130_fd_sc_hs__fill_2 FILLER_122_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_122_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_122_307 ();
 sky130_fd_sc_hs__fill_4 FILLER_122_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_122_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_122_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_122_336 ();
 sky130_fd_sc_hs__fill_1 FILLER_122_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_122_358 ();
 sky130_fd_sc_hs__fill_8 FILLER_122_366 ();
 sky130_fd_sc_hs__fill_2 FILLER_122_374 ();
 sky130_fd_sc_hs__fill_1 FILLER_122_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_122_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_122_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_122_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_122_402 ();
 sky130_fd_sc_hs__fill_1 FILLER_122_410 ();
 sky130_fd_sc_hs__fill_2 FILLER_122_422 ();
 sky130_fd_sc_hs__fill_2 FILLER_122_433 ();
 sky130_fd_sc_hs__fill_4 FILLER_122_460 ();
 sky130_fd_sc_hs__fill_1 FILLER_122_464 ();
 sky130_fd_sc_hs__fill_4 FILLER_122_488 ();
 sky130_fd_sc_hs__fill_1 FILLER_122_492 ();
 sky130_fd_sc_hs__fill_2 FILLER_122_514 ();
 sky130_fd_sc_hs__fill_1 FILLER_122_539 ();
 sky130_fd_sc_hs__fill_4 FILLER_123_0 ();
 sky130_fd_sc_hs__fill_1 FILLER_123_4 ();
 sky130_fd_sc_hs__fill_8 FILLER_123_13 ();
 sky130_fd_sc_hs__fill_8 FILLER_123_21 ();
 sky130_fd_sc_hs__fill_8 FILLER_123_29 ();
 sky130_fd_sc_hs__fill_8 FILLER_123_37 ();
 sky130_fd_sc_hs__fill_8 FILLER_123_45 ();
 sky130_fd_sc_hs__fill_4 FILLER_123_53 ();
 sky130_fd_sc_hs__fill_1 FILLER_123_57 ();
 sky130_fd_sc_hs__fill_8 FILLER_123_59 ();
 sky130_fd_sc_hs__fill_1 FILLER_123_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_123_85 ();
 sky130_fd_sc_hs__fill_4 FILLER_123_93 ();
 sky130_fd_sc_hs__fill_2 FILLER_123_97 ();
 sky130_fd_sc_hs__fill_1 FILLER_123_99 ();
 sky130_fd_sc_hs__fill_4 FILLER_123_117 ();
 sky130_fd_sc_hs__fill_1 FILLER_123_121 ();
 sky130_fd_sc_hs__fill_8 FILLER_123_128 ();
 sky130_fd_sc_hs__fill_4 FILLER_123_136 ();
 sky130_fd_sc_hs__fill_4 FILLER_123_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_123_175 ();
 sky130_fd_sc_hs__fill_2 FILLER_123_183 ();
 sky130_fd_sc_hs__fill_1 FILLER_123_185 ();
 sky130_fd_sc_hs__fill_8 FILLER_123_214 ();
 sky130_fd_sc_hs__fill_8 FILLER_123_222 ();
 sky130_fd_sc_hs__fill_2 FILLER_123_230 ();
 sky130_fd_sc_hs__fill_8 FILLER_123_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_123_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_123_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_123_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_123_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_123_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_123_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_123_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_123_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_123_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_123_307 ();
 sky130_fd_sc_hs__fill_2 FILLER_123_315 ();
 sky130_fd_sc_hs__fill_1 FILLER_123_317 ();
 sky130_fd_sc_hs__fill_2 FILLER_123_326 ();
 sky130_fd_sc_hs__fill_1 FILLER_123_328 ();
 sky130_fd_sc_hs__fill_4 FILLER_123_333 ();
 sky130_fd_sc_hs__fill_1 FILLER_123_337 ();
 sky130_fd_sc_hs__fill_4 FILLER_123_341 ();
 sky130_fd_sc_hs__fill_2 FILLER_123_345 ();
 sky130_fd_sc_hs__fill_1 FILLER_123_347 ();
 sky130_fd_sc_hs__fill_2 FILLER_123_349 ();
 sky130_fd_sc_hs__fill_1 FILLER_123_351 ();
 sky130_fd_sc_hs__fill_8 FILLER_123_355 ();
 sky130_fd_sc_hs__fill_4 FILLER_123_363 ();
 sky130_fd_sc_hs__fill_8 FILLER_123_379 ();
 sky130_fd_sc_hs__fill_2 FILLER_123_387 ();
 sky130_fd_sc_hs__fill_8 FILLER_123_395 ();
 sky130_fd_sc_hs__fill_2 FILLER_123_403 ();
 sky130_fd_sc_hs__fill_1 FILLER_123_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_123_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_123_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_123_423 ();
 sky130_fd_sc_hs__fill_4 FILLER_123_431 ();
 sky130_fd_sc_hs__fill_1 FILLER_123_435 ();
 sky130_fd_sc_hs__fill_8 FILLER_123_450 ();
 sky130_fd_sc_hs__fill_4 FILLER_123_458 ();
 sky130_fd_sc_hs__fill_2 FILLER_123_462 ();
 sky130_fd_sc_hs__fill_8 FILLER_123_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_123_473 ();
 sky130_fd_sc_hs__fill_2 FILLER_123_481 ();
 sky130_fd_sc_hs__fill_2 FILLER_123_523 ();
 sky130_fd_sc_hs__fill_1 FILLER_123_525 ();
 sky130_fd_sc_hs__fill_2 FILLER_123_537 ();
 sky130_fd_sc_hs__fill_1 FILLER_123_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_124_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_124_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_124_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_124_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_124_28 ();
 sky130_fd_sc_hs__fill_4 FILLER_124_30 ();
 sky130_fd_sc_hs__fill_2 FILLER_124_34 ();
 sky130_fd_sc_hs__fill_1 FILLER_124_39 ();
 sky130_fd_sc_hs__fill_4 FILLER_124_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_124_62 ();
 sky130_fd_sc_hs__fill_2 FILLER_124_70 ();
 sky130_fd_sc_hs__fill_1 FILLER_124_72 ();
 sky130_fd_sc_hs__fill_8 FILLER_124_76 ();
 sky130_fd_sc_hs__fill_2 FILLER_124_84 ();
 sky130_fd_sc_hs__fill_1 FILLER_124_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_124_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_124_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_124_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_124_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_124_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_124_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_124_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_124_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_124_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_124_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_124_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_124_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_124_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_124_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_124_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_124_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_124_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_124_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_124_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_124_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_124_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_124_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_124_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_124_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_124_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_124_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_124_278 ();
 sky130_fd_sc_hs__fill_4 FILLER_124_286 ();
 sky130_fd_sc_hs__fill_1 FILLER_124_290 ();
 sky130_fd_sc_hs__fill_8 FILLER_124_304 ();
 sky130_fd_sc_hs__fill_4 FILLER_124_312 ();
 sky130_fd_sc_hs__fill_2 FILLER_124_316 ();
 sky130_fd_sc_hs__fill_1 FILLER_124_318 ();
 sky130_fd_sc_hs__fill_1 FILLER_124_326 ();
 sky130_fd_sc_hs__fill_8 FILLER_124_333 ();
 sky130_fd_sc_hs__fill_8 FILLER_124_341 ();
 sky130_fd_sc_hs__fill_2 FILLER_124_349 ();
 sky130_fd_sc_hs__fill_2 FILLER_124_354 ();
 sky130_fd_sc_hs__fill_1 FILLER_124_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_124_378 ();
 sky130_fd_sc_hs__fill_2 FILLER_124_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_124_410 ();
 sky130_fd_sc_hs__fill_1 FILLER_124_418 ();
 sky130_fd_sc_hs__fill_1 FILLER_124_423 ();
 sky130_fd_sc_hs__fill_4 FILLER_124_429 ();
 sky130_fd_sc_hs__fill_2 FILLER_124_433 ();
 sky130_fd_sc_hs__fill_8 FILLER_124_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_124_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_124_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_124_460 ();
 sky130_fd_sc_hs__fill_4 FILLER_124_468 ();
 sky130_fd_sc_hs__fill_2 FILLER_124_472 ();
 sky130_fd_sc_hs__fill_1 FILLER_124_474 ();
 sky130_fd_sc_hs__fill_4 FILLER_124_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_124_506 ();
 sky130_fd_sc_hs__fill_1 FILLER_124_520 ();
 sky130_fd_sc_hs__fill_8 FILLER_125_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_125_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_125_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_125_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_125_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_125_49 ();
 sky130_fd_sc_hs__fill_1 FILLER_125_57 ();
 sky130_fd_sc_hs__fill_8 FILLER_125_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_125_67 ();
 sky130_fd_sc_hs__fill_4 FILLER_125_75 ();
 sky130_fd_sc_hs__fill_1 FILLER_125_79 ();
 sky130_fd_sc_hs__fill_8 FILLER_125_84 ();
 sky130_fd_sc_hs__fill_4 FILLER_125_92 ();
 sky130_fd_sc_hs__fill_1 FILLER_125_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_125_101 ();
 sky130_fd_sc_hs__fill_4 FILLER_125_109 ();
 sky130_fd_sc_hs__fill_2 FILLER_125_113 ();
 sky130_fd_sc_hs__fill_1 FILLER_125_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_125_117 ();
 sky130_fd_sc_hs__fill_2 FILLER_125_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_125_147 ();
 sky130_fd_sc_hs__fill_8 FILLER_125_155 ();
 sky130_fd_sc_hs__fill_8 FILLER_125_163 ();
 sky130_fd_sc_hs__fill_2 FILLER_125_171 ();
 sky130_fd_sc_hs__fill_1 FILLER_125_173 ();
 sky130_fd_sc_hs__fill_2 FILLER_125_198 ();
 sky130_fd_sc_hs__fill_8 FILLER_125_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_125_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_125_220 ();
 sky130_fd_sc_hs__fill_4 FILLER_125_228 ();
 sky130_fd_sc_hs__fill_2 FILLER_125_233 ();
 sky130_fd_sc_hs__fill_1 FILLER_125_235 ();
 sky130_fd_sc_hs__fill_8 FILLER_125_266 ();
 sky130_fd_sc_hs__fill_1 FILLER_125_277 ();
 sky130_fd_sc_hs__fill_4 FILLER_125_285 ();
 sky130_fd_sc_hs__fill_1 FILLER_125_289 ();
 sky130_fd_sc_hs__fill_1 FILLER_125_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_125_303 ();
 sky130_fd_sc_hs__fill_4 FILLER_125_311 ();
 sky130_fd_sc_hs__fill_2 FILLER_125_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_125_338 ();
 sky130_fd_sc_hs__fill_2 FILLER_125_346 ();
 sky130_fd_sc_hs__fill_1 FILLER_125_349 ();
 sky130_fd_sc_hs__fill_2 FILLER_125_378 ();
 sky130_fd_sc_hs__fill_2 FILLER_125_388 ();
 sky130_fd_sc_hs__fill_4 FILLER_125_395 ();
 sky130_fd_sc_hs__fill_2 FILLER_125_399 ();
 sky130_fd_sc_hs__fill_2 FILLER_125_419 ();
 sky130_fd_sc_hs__fill_8 FILLER_125_427 ();
 sky130_fd_sc_hs__fill_8 FILLER_125_435 ();
 sky130_fd_sc_hs__fill_8 FILLER_125_443 ();
 sky130_fd_sc_hs__fill_8 FILLER_125_451 ();
 sky130_fd_sc_hs__fill_4 FILLER_125_459 ();
 sky130_fd_sc_hs__fill_1 FILLER_125_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_125_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_125_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_125_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_125_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_125_497 ();
 sky130_fd_sc_hs__fill_4 FILLER_125_505 ();
 sky130_fd_sc_hs__fill_2 FILLER_125_509 ();
 sky130_fd_sc_hs__fill_1 FILLER_125_511 ();
 sky130_fd_sc_hs__fill_1 FILLER_125_517 ();
 sky130_fd_sc_hs__fill_8 FILLER_125_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_125_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_125_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_126_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_126_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_126_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_126_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_126_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_126_30 ();
 sky130_fd_sc_hs__fill_4 FILLER_126_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_126_46 ();
 sky130_fd_sc_hs__fill_1 FILLER_126_54 ();
 sky130_fd_sc_hs__fill_2 FILLER_126_77 ();
 sky130_fd_sc_hs__fill_1 FILLER_126_82 ();
 sky130_fd_sc_hs__fill_2 FILLER_126_106 ();
 sky130_fd_sc_hs__fill_1 FILLER_126_108 ();
 sky130_fd_sc_hs__fill_8 FILLER_126_112 ();
 sky130_fd_sc_hs__fill_4 FILLER_126_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_126_135 ();
 sky130_fd_sc_hs__fill_2 FILLER_126_143 ();
 sky130_fd_sc_hs__fill_1 FILLER_126_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_126_176 ();
 sky130_fd_sc_hs__fill_8 FILLER_126_184 ();
 sky130_fd_sc_hs__fill_8 FILLER_126_192 ();
 sky130_fd_sc_hs__fill_2 FILLER_126_200 ();
 sky130_fd_sc_hs__fill_1 FILLER_126_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_126_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_126_212 ();
 sky130_fd_sc_hs__fill_4 FILLER_126_220 ();
 sky130_fd_sc_hs__fill_1 FILLER_126_224 ();
 sky130_fd_sc_hs__fill_4 FILLER_126_239 ();
 sky130_fd_sc_hs__fill_8 FILLER_126_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_126_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_126_262 ();
 sky130_fd_sc_hs__fill_4 FILLER_126_270 ();
 sky130_fd_sc_hs__fill_2 FILLER_126_274 ();
 sky130_fd_sc_hs__fill_2 FILLER_126_285 ();
 sky130_fd_sc_hs__fill_1 FILLER_126_287 ();
 sky130_fd_sc_hs__fill_2 FILLER_126_291 ();
 sky130_fd_sc_hs__fill_1 FILLER_126_293 ();
 sky130_fd_sc_hs__fill_1 FILLER_126_297 ();
 sky130_fd_sc_hs__fill_8 FILLER_126_304 ();
 sky130_fd_sc_hs__fill_4 FILLER_126_312 ();
 sky130_fd_sc_hs__fill_2 FILLER_126_316 ();
 sky130_fd_sc_hs__fill_1 FILLER_126_318 ();
 sky130_fd_sc_hs__fill_2 FILLER_126_320 ();
 sky130_fd_sc_hs__fill_1 FILLER_126_322 ();
 sky130_fd_sc_hs__fill_8 FILLER_126_335 ();
 sky130_fd_sc_hs__fill_4 FILLER_126_343 ();
 sky130_fd_sc_hs__fill_2 FILLER_126_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_126_355 ();
 sky130_fd_sc_hs__fill_2 FILLER_126_363 ();
 sky130_fd_sc_hs__fill_1 FILLER_126_378 ();
 sky130_fd_sc_hs__fill_4 FILLER_126_408 ();
 sky130_fd_sc_hs__fill_2 FILLER_126_412 ();
 sky130_fd_sc_hs__fill_8 FILLER_126_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_126_434 ();
 sky130_fd_sc_hs__fill_2 FILLER_126_436 ();
 sky130_fd_sc_hs__fill_1 FILLER_126_438 ();
 sky130_fd_sc_hs__fill_8 FILLER_126_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_126_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_126_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_126_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_126_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_126_492 ();
 sky130_fd_sc_hs__fill_4 FILLER_126_494 ();
 sky130_fd_sc_hs__fill_2 FILLER_126_498 ();
 sky130_fd_sc_hs__fill_8 FILLER_126_508 ();
 sky130_fd_sc_hs__fill_8 FILLER_126_516 ();
 sky130_fd_sc_hs__fill_8 FILLER_126_524 ();
 sky130_fd_sc_hs__fill_8 FILLER_127_0 ();
 sky130_fd_sc_hs__fill_4 FILLER_127_8 ();
 sky130_fd_sc_hs__fill_1 FILLER_127_12 ();
 sky130_fd_sc_hs__fill_8 FILLER_127_21 ();
 sky130_fd_sc_hs__fill_8 FILLER_127_29 ();
 sky130_fd_sc_hs__fill_8 FILLER_127_37 ();
 sky130_fd_sc_hs__fill_8 FILLER_127_45 ();
 sky130_fd_sc_hs__fill_4 FILLER_127_53 ();
 sky130_fd_sc_hs__fill_1 FILLER_127_57 ();
 sky130_fd_sc_hs__fill_4 FILLER_127_59 ();
 sky130_fd_sc_hs__fill_2 FILLER_127_63 ();
 sky130_fd_sc_hs__fill_2 FILLER_127_95 ();
 sky130_fd_sc_hs__fill_1 FILLER_127_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_127_138 ();
 sky130_fd_sc_hs__fill_8 FILLER_127_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_127_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_127_162 ();
 sky130_fd_sc_hs__fill_4 FILLER_127_170 ();
 sky130_fd_sc_hs__fill_4 FILLER_127_181 ();
 sky130_fd_sc_hs__fill_2 FILLER_127_193 ();
 sky130_fd_sc_hs__fill_8 FILLER_127_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_127_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_127_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_127_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_127_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_127_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_127_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_127_273 ();
 sky130_fd_sc_hs__fill_2 FILLER_127_291 ();
 sky130_fd_sc_hs__fill_1 FILLER_127_293 ();
 sky130_fd_sc_hs__fill_8 FILLER_127_311 ();
 sky130_fd_sc_hs__fill_8 FILLER_127_319 ();
 sky130_fd_sc_hs__fill_8 FILLER_127_327 ();
 sky130_fd_sc_hs__fill_4 FILLER_127_335 ();
 sky130_fd_sc_hs__fill_2 FILLER_127_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_127_341 ();
 sky130_fd_sc_hs__fill_2 FILLER_127_345 ();
 sky130_fd_sc_hs__fill_1 FILLER_127_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_127_349 ();
 sky130_fd_sc_hs__fill_4 FILLER_127_357 ();
 sky130_fd_sc_hs__fill_1 FILLER_127_361 ();
 sky130_fd_sc_hs__fill_8 FILLER_127_388 ();
 sky130_fd_sc_hs__fill_8 FILLER_127_396 ();
 sky130_fd_sc_hs__fill_2 FILLER_127_404 ();
 sky130_fd_sc_hs__fill_1 FILLER_127_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_127_424 ();
 sky130_fd_sc_hs__fill_8 FILLER_127_432 ();
 sky130_fd_sc_hs__fill_8 FILLER_127_452 ();
 sky130_fd_sc_hs__fill_4 FILLER_127_460 ();
 sky130_fd_sc_hs__fill_4 FILLER_127_465 ();
 sky130_fd_sc_hs__fill_1 FILLER_127_469 ();
 sky130_fd_sc_hs__fill_8 FILLER_127_487 ();
 sky130_fd_sc_hs__fill_8 FILLER_127_495 ();
 sky130_fd_sc_hs__fill_8 FILLER_127_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_127_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_127_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_128_0 ();
 sky130_fd_sc_hs__fill_4 FILLER_128_8 ();
 sky130_fd_sc_hs__fill_2 FILLER_128_12 ();
 sky130_fd_sc_hs__fill_4 FILLER_128_22 ();
 sky130_fd_sc_hs__fill_2 FILLER_128_26 ();
 sky130_fd_sc_hs__fill_1 FILLER_128_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_128_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_128_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_128_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_128_88 ();
 sky130_fd_sc_hs__fill_2 FILLER_128_106 ();
 sky130_fd_sc_hs__fill_8 FILLER_128_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_128_144 ();
 sky130_fd_sc_hs__fill_4 FILLER_128_146 ();
 sky130_fd_sc_hs__fill_1 FILLER_128_150 ();
 sky130_fd_sc_hs__fill_8 FILLER_128_174 ();
 sky130_fd_sc_hs__fill_2 FILLER_128_182 ();
 sky130_fd_sc_hs__fill_8 FILLER_128_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_128_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_128_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_128_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_128_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_128_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_128_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_128_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_128_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_128_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_128_269 ();
 sky130_fd_sc_hs__fill_1 FILLER_128_277 ();
 sky130_fd_sc_hs__fill_1 FILLER_128_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_128_304 ();
 sky130_fd_sc_hs__fill_4 FILLER_128_312 ();
 sky130_fd_sc_hs__fill_2 FILLER_128_316 ();
 sky130_fd_sc_hs__fill_1 FILLER_128_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_128_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_128_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_128_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_128_344 ();
 sky130_fd_sc_hs__fill_4 FILLER_128_352 ();
 sky130_fd_sc_hs__fill_1 FILLER_128_356 ();
 sky130_fd_sc_hs__fill_8 FILLER_128_365 ();
 sky130_fd_sc_hs__fill_4 FILLER_128_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_128_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_128_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_128_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_128_402 ();
 sky130_fd_sc_hs__fill_2 FILLER_128_410 ();
 sky130_fd_sc_hs__fill_4 FILLER_128_436 ();
 sky130_fd_sc_hs__fill_1 FILLER_128_452 ();
 sky130_fd_sc_hs__fill_4 FILLER_128_488 ();
 sky130_fd_sc_hs__fill_1 FILLER_128_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_128_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_128_502 ();
 sky130_fd_sc_hs__fill_1 FILLER_128_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_129_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_129_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_129_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_129_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_129_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_129_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_129_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_129_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_129_67 ();
 sky130_fd_sc_hs__fill_4 FILLER_129_75 ();
 sky130_fd_sc_hs__fill_2 FILLER_129_79 ();
 sky130_fd_sc_hs__fill_1 FILLER_129_81 ();
 sky130_fd_sc_hs__fill_8 FILLER_129_90 ();
 sky130_fd_sc_hs__fill_8 FILLER_129_126 ();
 sky130_fd_sc_hs__fill_2 FILLER_129_134 ();
 sky130_fd_sc_hs__fill_1 FILLER_129_136 ();
 sky130_fd_sc_hs__fill_8 FILLER_129_162 ();
 sky130_fd_sc_hs__fill_1 FILLER_129_170 ();
 sky130_fd_sc_hs__fill_1 FILLER_129_175 ();
 sky130_fd_sc_hs__fill_1 FILLER_129_191 ();
 sky130_fd_sc_hs__fill_2 FILLER_129_200 ();
 sky130_fd_sc_hs__fill_1 FILLER_129_202 ();
 sky130_fd_sc_hs__fill_2 FILLER_129_206 ();
 sky130_fd_sc_hs__fill_4 FILLER_129_227 ();
 sky130_fd_sc_hs__fill_1 FILLER_129_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_129_233 ();
 sky130_fd_sc_hs__fill_4 FILLER_129_241 ();
 sky130_fd_sc_hs__fill_1 FILLER_129_245 ();
 sky130_fd_sc_hs__fill_8 FILLER_129_272 ();
 sky130_fd_sc_hs__fill_4 FILLER_129_280 ();
 sky130_fd_sc_hs__fill_1 FILLER_129_284 ();
 sky130_fd_sc_hs__fill_1 FILLER_129_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_129_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_129_302 ();
 sky130_fd_sc_hs__fill_8 FILLER_129_310 ();
 sky130_fd_sc_hs__fill_8 FILLER_129_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_129_326 ();
 sky130_fd_sc_hs__fill_8 FILLER_129_334 ();
 sky130_fd_sc_hs__fill_4 FILLER_129_342 ();
 sky130_fd_sc_hs__fill_2 FILLER_129_346 ();
 sky130_fd_sc_hs__fill_8 FILLER_129_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_129_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_129_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_129_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_129_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_129_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_129_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_129_405 ();
 sky130_fd_sc_hs__fill_1 FILLER_129_407 ();
 sky130_fd_sc_hs__fill_4 FILLER_129_420 ();
 sky130_fd_sc_hs__fill_2 FILLER_129_424 ();
 sky130_fd_sc_hs__fill_1 FILLER_129_426 ();
 sky130_fd_sc_hs__fill_8 FILLER_129_435 ();
 sky130_fd_sc_hs__fill_8 FILLER_129_443 ();
 sky130_fd_sc_hs__fill_8 FILLER_129_451 ();
 sky130_fd_sc_hs__fill_4 FILLER_129_459 ();
 sky130_fd_sc_hs__fill_1 FILLER_129_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_129_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_129_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_129_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_129_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_129_497 ();
 sky130_fd_sc_hs__fill_4 FILLER_129_505 ();
 sky130_fd_sc_hs__fill_2 FILLER_129_509 ();
 sky130_fd_sc_hs__fill_2 FILLER_129_520 ();
 sky130_fd_sc_hs__fill_2 FILLER_129_523 ();
 sky130_fd_sc_hs__fill_1 FILLER_129_525 ();
 sky130_fd_sc_hs__fill_2 FILLER_129_537 ();
 sky130_fd_sc_hs__fill_1 FILLER_129_539 ();
 sky130_fd_sc_hs__fill_4 FILLER_130_0 ();
 sky130_fd_sc_hs__fill_1 FILLER_130_4 ();
 sky130_fd_sc_hs__fill_8 FILLER_130_13 ();
 sky130_fd_sc_hs__fill_8 FILLER_130_21 ();
 sky130_fd_sc_hs__fill_8 FILLER_130_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_130_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_130_46 ();
 sky130_fd_sc_hs__fill_2 FILLER_130_54 ();
 sky130_fd_sc_hs__fill_2 FILLER_130_67 ();
 sky130_fd_sc_hs__fill_4 FILLER_130_73 ();
 sky130_fd_sc_hs__fill_1 FILLER_130_77 ();
 sky130_fd_sc_hs__fill_8 FILLER_130_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_130_96 ();
 sky130_fd_sc_hs__fill_2 FILLER_130_104 ();
 sky130_fd_sc_hs__fill_2 FILLER_130_109 ();
 sky130_fd_sc_hs__fill_1 FILLER_130_111 ();
 sky130_fd_sc_hs__fill_8 FILLER_130_116 ();
 sky130_fd_sc_hs__fill_8 FILLER_130_124 ();
 sky130_fd_sc_hs__fill_8 FILLER_130_132 ();
 sky130_fd_sc_hs__fill_8 FILLER_130_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_130_190 ();
 sky130_fd_sc_hs__fill_4 FILLER_130_198 ();
 sky130_fd_sc_hs__fill_1 FILLER_130_202 ();
 sky130_fd_sc_hs__fill_2 FILLER_130_204 ();
 sky130_fd_sc_hs__fill_1 FILLER_130_206 ();
 sky130_fd_sc_hs__fill_8 FILLER_130_226 ();
 sky130_fd_sc_hs__fill_2 FILLER_130_234 ();
 sky130_fd_sc_hs__fill_4 FILLER_130_239 ();
 sky130_fd_sc_hs__fill_8 FILLER_130_250 ();
 sky130_fd_sc_hs__fill_2 FILLER_130_258 ();
 sky130_fd_sc_hs__fill_1 FILLER_130_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_130_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_130_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_130_278 ();
 sky130_fd_sc_hs__fill_1 FILLER_130_286 ();
 sky130_fd_sc_hs__fill_4 FILLER_130_296 ();
 sky130_fd_sc_hs__fill_2 FILLER_130_312 ();
 sky130_fd_sc_hs__fill_1 FILLER_130_314 ();
 sky130_fd_sc_hs__fill_1 FILLER_130_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_130_326 ();
 sky130_fd_sc_hs__fill_2 FILLER_130_334 ();
 sky130_fd_sc_hs__fill_4 FILLER_130_345 ();
 sky130_fd_sc_hs__fill_8 FILLER_130_354 ();
 sky130_fd_sc_hs__fill_8 FILLER_130_362 ();
 sky130_fd_sc_hs__fill_4 FILLER_130_370 ();
 sky130_fd_sc_hs__fill_2 FILLER_130_374 ();
 sky130_fd_sc_hs__fill_1 FILLER_130_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_130_378 ();
 sky130_fd_sc_hs__fill_2 FILLER_130_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_130_395 ();
 sky130_fd_sc_hs__fill_8 FILLER_130_403 ();
 sky130_fd_sc_hs__fill_8 FILLER_130_411 ();
 sky130_fd_sc_hs__fill_4 FILLER_130_419 ();
 sky130_fd_sc_hs__fill_2 FILLER_130_423 ();
 sky130_fd_sc_hs__fill_1 FILLER_130_425 ();
 sky130_fd_sc_hs__fill_8 FILLER_130_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_130_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_130_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_130_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_130_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_130_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_130_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_130_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_130_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_130_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_130_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_130_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_130_526 ();
 sky130_fd_sc_hs__fill_4 FILLER_130_534 ();
 sky130_fd_sc_hs__fill_2 FILLER_130_538 ();
 sky130_fd_sc_hs__fill_8 FILLER_131_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_131_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_131_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_131_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_131_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_131_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_131_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_131_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_131_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_131_87 ();
 sky130_fd_sc_hs__fill_8 FILLER_131_95 ();
 sky130_fd_sc_hs__fill_8 FILLER_131_103 ();
 sky130_fd_sc_hs__fill_4 FILLER_131_111 ();
 sky130_fd_sc_hs__fill_1 FILLER_131_115 ();
 sky130_fd_sc_hs__fill_4 FILLER_131_117 ();
 sky130_fd_sc_hs__fill_2 FILLER_131_121 ();
 sky130_fd_sc_hs__fill_4 FILLER_131_126 ();
 sky130_fd_sc_hs__fill_2 FILLER_131_130 ();
 sky130_fd_sc_hs__fill_1 FILLER_131_132 ();
 sky130_fd_sc_hs__fill_8 FILLER_131_145 ();
 sky130_fd_sc_hs__fill_8 FILLER_131_153 ();
 sky130_fd_sc_hs__fill_8 FILLER_131_161 ();
 sky130_fd_sc_hs__fill_4 FILLER_131_169 ();
 sky130_fd_sc_hs__fill_1 FILLER_131_173 ();
 sky130_fd_sc_hs__fill_4 FILLER_131_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_131_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_131_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_131_220 ();
 sky130_fd_sc_hs__fill_4 FILLER_131_228 ();
 sky130_fd_sc_hs__fill_2 FILLER_131_233 ();
 sky130_fd_sc_hs__fill_1 FILLER_131_235 ();
 sky130_fd_sc_hs__fill_2 FILLER_131_239 ();
 sky130_fd_sc_hs__fill_1 FILLER_131_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_131_246 ();
 sky130_fd_sc_hs__fill_8 FILLER_131_254 ();
 sky130_fd_sc_hs__fill_8 FILLER_131_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_131_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_131_278 ();
 sky130_fd_sc_hs__fill_4 FILLER_131_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_131_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_131_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_131_307 ();
 sky130_fd_sc_hs__fill_2 FILLER_131_315 ();
 sky130_fd_sc_hs__fill_1 FILLER_131_317 ();
 sky130_fd_sc_hs__fill_8 FILLER_131_325 ();
 sky130_fd_sc_hs__fill_4 FILLER_131_333 ();
 sky130_fd_sc_hs__fill_8 FILLER_131_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_131_357 ();
 sky130_fd_sc_hs__fill_1 FILLER_131_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_131_387 ();
 sky130_fd_sc_hs__fill_8 FILLER_131_395 ();
 sky130_fd_sc_hs__fill_2 FILLER_131_403 ();
 sky130_fd_sc_hs__fill_1 FILLER_131_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_131_416 ();
 sky130_fd_sc_hs__fill_8 FILLER_131_424 ();
 sky130_fd_sc_hs__fill_8 FILLER_131_432 ();
 sky130_fd_sc_hs__fill_8 FILLER_131_440 ();
 sky130_fd_sc_hs__fill_8 FILLER_131_448 ();
 sky130_fd_sc_hs__fill_1 FILLER_131_456 ();
 sky130_fd_sc_hs__fill_8 FILLER_131_465 ();
 sky130_fd_sc_hs__fill_2 FILLER_131_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_131_498 ();
 sky130_fd_sc_hs__fill_8 FILLER_131_523 ();
 sky130_fd_sc_hs__fill_1 FILLER_131_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_132_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_132_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_132_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_132_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_132_28 ();
 sky130_fd_sc_hs__fill_4 FILLER_132_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_132_51 ();
 sky130_fd_sc_hs__fill_8 FILLER_132_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_132_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_132_75 ();
 sky130_fd_sc_hs__fill_4 FILLER_132_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_132_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_132_126 ();
 sky130_fd_sc_hs__fill_4 FILLER_132_134 ();
 sky130_fd_sc_hs__fill_1 FILLER_132_138 ();
 sky130_fd_sc_hs__fill_8 FILLER_132_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_132_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_132_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_132_170 ();
 sky130_fd_sc_hs__fill_4 FILLER_132_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_132_204 ();
 sky130_fd_sc_hs__fill_2 FILLER_132_212 ();
 sky130_fd_sc_hs__fill_1 FILLER_132_214 ();
 sky130_fd_sc_hs__fill_8 FILLER_132_218 ();
 sky130_fd_sc_hs__fill_2 FILLER_132_226 ();
 sky130_fd_sc_hs__fill_1 FILLER_132_228 ();
 sky130_fd_sc_hs__fill_1 FILLER_132_243 ();
 sky130_fd_sc_hs__fill_8 FILLER_132_249 ();
 sky130_fd_sc_hs__fill_4 FILLER_132_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_132_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_132_283 ();
 sky130_fd_sc_hs__fill_8 FILLER_132_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_132_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_132_307 ();
 sky130_fd_sc_hs__fill_4 FILLER_132_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_132_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_132_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_132_339 ();
 sky130_fd_sc_hs__fill_8 FILLER_132_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_132_355 ();
 sky130_fd_sc_hs__fill_8 FILLER_132_363 ();
 sky130_fd_sc_hs__fill_4 FILLER_132_371 ();
 sky130_fd_sc_hs__fill_2 FILLER_132_375 ();
 sky130_fd_sc_hs__fill_8 FILLER_132_378 ();
 sky130_fd_sc_hs__fill_4 FILLER_132_386 ();
 sky130_fd_sc_hs__fill_2 FILLER_132_390 ();
 sky130_fd_sc_hs__fill_1 FILLER_132_392 ();
 sky130_fd_sc_hs__fill_4 FILLER_132_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_132_436 ();
 sky130_fd_sc_hs__fill_2 FILLER_132_457 ();
 sky130_fd_sc_hs__fill_1 FILLER_132_459 ();
 sky130_fd_sc_hs__fill_2 FILLER_132_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_132_516 ();
 sky130_fd_sc_hs__fill_8 FILLER_132_524 ();
 sky130_fd_sc_hs__fill_8 FILLER_133_0 ();
 sky130_fd_sc_hs__fill_2 FILLER_133_8 ();
 sky130_fd_sc_hs__fill_1 FILLER_133_10 ();
 sky130_fd_sc_hs__fill_8 FILLER_133_27 ();
 sky130_fd_sc_hs__fill_1 FILLER_133_35 ();
 sky130_fd_sc_hs__fill_1 FILLER_133_57 ();
 sky130_fd_sc_hs__fill_8 FILLER_133_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_133_67 ();
 sky130_fd_sc_hs__fill_4 FILLER_133_75 ();
 sky130_fd_sc_hs__fill_4 FILLER_133_87 ();
 sky130_fd_sc_hs__fill_2 FILLER_133_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_133_101 ();
 sky130_fd_sc_hs__fill_4 FILLER_133_109 ();
 sky130_fd_sc_hs__fill_2 FILLER_133_113 ();
 sky130_fd_sc_hs__fill_1 FILLER_133_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_133_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_133_125 ();
 sky130_fd_sc_hs__fill_1 FILLER_133_173 ();
 sky130_fd_sc_hs__fill_2 FILLER_133_181 ();
 sky130_fd_sc_hs__fill_1 FILLER_133_187 ();
 sky130_fd_sc_hs__fill_8 FILLER_133_192 ();
 sky130_fd_sc_hs__fill_8 FILLER_133_200 ();
 sky130_fd_sc_hs__fill_2 FILLER_133_208 ();
 sky130_fd_sc_hs__fill_1 FILLER_133_210 ();
 sky130_fd_sc_hs__fill_4 FILLER_133_233 ();
 sky130_fd_sc_hs__fill_1 FILLER_133_237 ();
 sky130_fd_sc_hs__fill_8 FILLER_133_256 ();
 sky130_fd_sc_hs__fill_2 FILLER_133_270 ();
 sky130_fd_sc_hs__fill_1 FILLER_133_272 ();
 sky130_fd_sc_hs__fill_8 FILLER_133_277 ();
 sky130_fd_sc_hs__fill_4 FILLER_133_285 ();
 sky130_fd_sc_hs__fill_1 FILLER_133_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_133_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_133_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_133_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_133_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_133_323 ();
 sky130_fd_sc_hs__fill_4 FILLER_133_331 ();
 sky130_fd_sc_hs__fill_2 FILLER_133_335 ();
 sky130_fd_sc_hs__fill_8 FILLER_133_340 ();
 sky130_fd_sc_hs__fill_8 FILLER_133_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_133_357 ();
 sky130_fd_sc_hs__fill_1 FILLER_133_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_133_369 ();
 sky130_fd_sc_hs__fill_8 FILLER_133_377 ();
 sky130_fd_sc_hs__fill_8 FILLER_133_385 ();
 sky130_fd_sc_hs__fill_1 FILLER_133_393 ();
 sky130_fd_sc_hs__fill_8 FILLER_133_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_133_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_133_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_133_431 ();
 sky130_fd_sc_hs__fill_4 FILLER_133_439 ();
 sky130_fd_sc_hs__fill_2 FILLER_133_443 ();
 sky130_fd_sc_hs__fill_1 FILLER_133_445 ();
 sky130_fd_sc_hs__fill_8 FILLER_133_450 ();
 sky130_fd_sc_hs__fill_4 FILLER_133_458 ();
 sky130_fd_sc_hs__fill_2 FILLER_133_462 ();
 sky130_fd_sc_hs__fill_8 FILLER_133_465 ();
 sky130_fd_sc_hs__fill_4 FILLER_133_473 ();
 sky130_fd_sc_hs__fill_2 FILLER_133_477 ();
 sky130_fd_sc_hs__fill_1 FILLER_133_479 ();
 sky130_fd_sc_hs__fill_2 FILLER_133_500 ();
 sky130_fd_sc_hs__fill_8 FILLER_133_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_133_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_133_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_134_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_134_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_134_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_134_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_134_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_134_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_134_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_134_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_134_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_134_62 ();
 sky130_fd_sc_hs__fill_4 FILLER_134_70 ();
 sky130_fd_sc_hs__fill_2 FILLER_134_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_134_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_134_125 ();
 sky130_fd_sc_hs__fill_4 FILLER_134_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_134_146 ();
 sky130_fd_sc_hs__fill_4 FILLER_134_154 ();
 sky130_fd_sc_hs__fill_2 FILLER_134_158 ();
 sky130_fd_sc_hs__fill_1 FILLER_134_160 ();
 sky130_fd_sc_hs__fill_8 FILLER_134_169 ();
 sky130_fd_sc_hs__fill_8 FILLER_134_177 ();
 sky130_fd_sc_hs__fill_8 FILLER_134_185 ();
 sky130_fd_sc_hs__fill_8 FILLER_134_193 ();
 sky130_fd_sc_hs__fill_2 FILLER_134_201 ();
 sky130_fd_sc_hs__fill_8 FILLER_134_204 ();
 sky130_fd_sc_hs__fill_1 FILLER_134_212 ();
 sky130_fd_sc_hs__fill_2 FILLER_134_236 ();
 sky130_fd_sc_hs__fill_1 FILLER_134_238 ();
 sky130_fd_sc_hs__fill_2 FILLER_134_246 ();
 sky130_fd_sc_hs__fill_1 FILLER_134_248 ();
 sky130_fd_sc_hs__fill_8 FILLER_134_278 ();
 sky130_fd_sc_hs__fill_1 FILLER_134_286 ();
 sky130_fd_sc_hs__fill_4 FILLER_134_299 ();
 sky130_fd_sc_hs__fill_2 FILLER_134_303 ();
 sky130_fd_sc_hs__fill_1 FILLER_134_305 ();
 sky130_fd_sc_hs__fill_1 FILLER_134_320 ();
 sky130_fd_sc_hs__fill_1 FILLER_134_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_134_385 ();
 sky130_fd_sc_hs__fill_8 FILLER_134_393 ();
 sky130_fd_sc_hs__fill_8 FILLER_134_401 ();
 sky130_fd_sc_hs__fill_4 FILLER_134_409 ();
 sky130_fd_sc_hs__fill_2 FILLER_134_413 ();
 sky130_fd_sc_hs__fill_4 FILLER_134_431 ();
 sky130_fd_sc_hs__fill_1 FILLER_134_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_134_462 ();
 sky130_fd_sc_hs__fill_8 FILLER_134_470 ();
 sky130_fd_sc_hs__fill_8 FILLER_134_478 ();
 sky130_fd_sc_hs__fill_4 FILLER_134_486 ();
 sky130_fd_sc_hs__fill_2 FILLER_134_490 ();
 sky130_fd_sc_hs__fill_1 FILLER_134_492 ();
 sky130_fd_sc_hs__fill_2 FILLER_134_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_134_519 ();
 sky130_fd_sc_hs__fill_8 FILLER_134_527 ();
 sky130_fd_sc_hs__fill_4 FILLER_134_535 ();
 sky130_fd_sc_hs__fill_1 FILLER_134_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_135_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_135_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_135_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_135_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_135_28 ();
 sky130_fd_sc_hs__fill_2 FILLER_135_37 ();
 sky130_fd_sc_hs__fill_1 FILLER_135_39 ();
 sky130_fd_sc_hs__fill_8 FILLER_135_47 ();
 sky130_fd_sc_hs__fill_2 FILLER_135_55 ();
 sky130_fd_sc_hs__fill_1 FILLER_135_57 ();
 sky130_fd_sc_hs__fill_8 FILLER_135_59 ();
 sky130_fd_sc_hs__fill_4 FILLER_135_67 ();
 sky130_fd_sc_hs__fill_2 FILLER_135_71 ();
 sky130_fd_sc_hs__fill_8 FILLER_135_94 ();
 sky130_fd_sc_hs__fill_8 FILLER_135_102 ();
 sky130_fd_sc_hs__fill_4 FILLER_135_110 ();
 sky130_fd_sc_hs__fill_2 FILLER_135_114 ();
 sky130_fd_sc_hs__fill_8 FILLER_135_117 ();
 sky130_fd_sc_hs__fill_2 FILLER_135_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_135_154 ();
 sky130_fd_sc_hs__fill_4 FILLER_135_169 ();
 sky130_fd_sc_hs__fill_1 FILLER_135_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_135_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_135_183 ();
 sky130_fd_sc_hs__fill_4 FILLER_135_191 ();
 sky130_fd_sc_hs__fill_2 FILLER_135_195 ();
 sky130_fd_sc_hs__fill_1 FILLER_135_197 ();
 sky130_fd_sc_hs__fill_8 FILLER_135_209 ();
 sky130_fd_sc_hs__fill_8 FILLER_135_217 ();
 sky130_fd_sc_hs__fill_4 FILLER_135_225 ();
 sky130_fd_sc_hs__fill_2 FILLER_135_229 ();
 sky130_fd_sc_hs__fill_1 FILLER_135_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_135_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_135_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_135_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_135_269 ();
 sky130_fd_sc_hs__fill_8 FILLER_135_277 ();
 sky130_fd_sc_hs__fill_4 FILLER_135_285 ();
 sky130_fd_sc_hs__fill_1 FILLER_135_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_135_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_135_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_135_307 ();
 sky130_fd_sc_hs__fill_4 FILLER_135_315 ();
 sky130_fd_sc_hs__fill_1 FILLER_135_319 ();
 sky130_fd_sc_hs__fill_8 FILLER_135_333 ();
 sky130_fd_sc_hs__fill_4 FILLER_135_341 ();
 sky130_fd_sc_hs__fill_2 FILLER_135_345 ();
 sky130_fd_sc_hs__fill_1 FILLER_135_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_135_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_135_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_135_365 ();
 sky130_fd_sc_hs__fill_1 FILLER_135_373 ();
 sky130_fd_sc_hs__fill_1 FILLER_135_380 ();
 sky130_fd_sc_hs__fill_8 FILLER_135_390 ();
 sky130_fd_sc_hs__fill_8 FILLER_135_398 ();
 sky130_fd_sc_hs__fill_8 FILLER_135_407 ();
 sky130_fd_sc_hs__fill_2 FILLER_135_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_135_430 ();
 sky130_fd_sc_hs__fill_8 FILLER_135_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_135_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_135_477 ();
 sky130_fd_sc_hs__fill_8 FILLER_135_485 ();
 sky130_fd_sc_hs__fill_2 FILLER_135_493 ();
 sky130_fd_sc_hs__fill_2 FILLER_135_501 ();
 sky130_fd_sc_hs__fill_2 FILLER_135_537 ();
 sky130_fd_sc_hs__fill_1 FILLER_135_539 ();
 sky130_fd_sc_hs__fill_4 FILLER_136_0 ();
 sky130_fd_sc_hs__fill_1 FILLER_136_4 ();
 sky130_fd_sc_hs__fill_8 FILLER_136_13 ();
 sky130_fd_sc_hs__fill_8 FILLER_136_21 ();
 sky130_fd_sc_hs__fill_8 FILLER_136_30 ();
 sky130_fd_sc_hs__fill_1 FILLER_136_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_136_65 ();
 sky130_fd_sc_hs__fill_2 FILLER_136_73 ();
 sky130_fd_sc_hs__fill_1 FILLER_136_75 ();
 sky130_fd_sc_hs__fill_1 FILLER_136_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_136_107 ();
 sky130_fd_sc_hs__fill_8 FILLER_136_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_136_123 ();
 sky130_fd_sc_hs__fill_2 FILLER_136_131 ();
 sky130_fd_sc_hs__fill_4 FILLER_136_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_136_176 ();
 sky130_fd_sc_hs__fill_4 FILLER_136_184 ();
 sky130_fd_sc_hs__fill_2 FILLER_136_188 ();
 sky130_fd_sc_hs__fill_1 FILLER_136_190 ();
 sky130_fd_sc_hs__fill_8 FILLER_136_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_136_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_136_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_136_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_136_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_136_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_136_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_136_260 ();
 sky130_fd_sc_hs__fill_4 FILLER_136_262 ();
 sky130_fd_sc_hs__fill_1 FILLER_136_266 ();
 sky130_fd_sc_hs__fill_8 FILLER_136_270 ();
 sky130_fd_sc_hs__fill_4 FILLER_136_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_136_288 ();
 sky130_fd_sc_hs__fill_8 FILLER_136_296 ();
 sky130_fd_sc_hs__fill_8 FILLER_136_304 ();
 sky130_fd_sc_hs__fill_4 FILLER_136_312 ();
 sky130_fd_sc_hs__fill_2 FILLER_136_316 ();
 sky130_fd_sc_hs__fill_1 FILLER_136_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_136_327 ();
 sky130_fd_sc_hs__fill_8 FILLER_136_335 ();
 sky130_fd_sc_hs__fill_8 FILLER_136_343 ();
 sky130_fd_sc_hs__fill_8 FILLER_136_351 ();
 sky130_fd_sc_hs__fill_8 FILLER_136_359 ();
 sky130_fd_sc_hs__fill_8 FILLER_136_367 ();
 sky130_fd_sc_hs__fill_2 FILLER_136_375 ();
 sky130_fd_sc_hs__fill_8 FILLER_136_390 ();
 sky130_fd_sc_hs__fill_1 FILLER_136_398 ();
 sky130_fd_sc_hs__fill_8 FILLER_136_404 ();
 sky130_fd_sc_hs__fill_4 FILLER_136_412 ();
 sky130_fd_sc_hs__fill_2 FILLER_136_416 ();
 sky130_fd_sc_hs__fill_1 FILLER_136_418 ();
 sky130_fd_sc_hs__fill_4 FILLER_136_430 ();
 sky130_fd_sc_hs__fill_1 FILLER_136_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_136_436 ();
 sky130_fd_sc_hs__fill_2 FILLER_136_444 ();
 sky130_fd_sc_hs__fill_4 FILLER_136_458 ();
 sky130_fd_sc_hs__fill_2 FILLER_136_462 ();
 sky130_fd_sc_hs__fill_8 FILLER_136_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_136_481 ();
 sky130_fd_sc_hs__fill_4 FILLER_136_489 ();
 sky130_fd_sc_hs__fill_4 FILLER_136_494 ();
 sky130_fd_sc_hs__fill_2 FILLER_136_498 ();
 sky130_fd_sc_hs__fill_2 FILLER_136_506 ();
 sky130_fd_sc_hs__fill_8 FILLER_137_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_137_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_137_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_137_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_137_32 ();
 sky130_fd_sc_hs__fill_4 FILLER_137_40 ();
 sky130_fd_sc_hs__fill_4 FILLER_137_53 ();
 sky130_fd_sc_hs__fill_1 FILLER_137_57 ();
 sky130_fd_sc_hs__fill_8 FILLER_137_59 ();
 sky130_fd_sc_hs__fill_4 FILLER_137_67 ();
 sky130_fd_sc_hs__fill_1 FILLER_137_71 ();
 sky130_fd_sc_hs__fill_2 FILLER_137_78 ();
 sky130_fd_sc_hs__fill_8 FILLER_137_105 ();
 sky130_fd_sc_hs__fill_2 FILLER_137_113 ();
 sky130_fd_sc_hs__fill_1 FILLER_137_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_137_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_137_146 ();
 sky130_fd_sc_hs__fill_4 FILLER_137_154 ();
 sky130_fd_sc_hs__fill_2 FILLER_137_158 ();
 sky130_fd_sc_hs__fill_1 FILLER_137_160 ();
 sky130_fd_sc_hs__fill_1 FILLER_137_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_137_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_137_183 ();
 sky130_fd_sc_hs__fill_1 FILLER_137_195 ();
 sky130_fd_sc_hs__fill_8 FILLER_137_208 ();
 sky130_fd_sc_hs__fill_8 FILLER_137_216 ();
 sky130_fd_sc_hs__fill_8 FILLER_137_224 ();
 sky130_fd_sc_hs__fill_8 FILLER_137_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_137_241 ();
 sky130_fd_sc_hs__fill_2 FILLER_137_249 ();
 sky130_fd_sc_hs__fill_1 FILLER_137_251 ();
 sky130_fd_sc_hs__fill_8 FILLER_137_271 ();
 sky130_fd_sc_hs__fill_8 FILLER_137_279 ();
 sky130_fd_sc_hs__fill_2 FILLER_137_287 ();
 sky130_fd_sc_hs__fill_1 FILLER_137_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_137_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_137_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_137_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_137_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_137_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_137_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_137_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_137_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_137_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_137_357 ();
 sky130_fd_sc_hs__fill_1 FILLER_137_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_137_389 ();
 sky130_fd_sc_hs__fill_2 FILLER_137_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_137_399 ();
 sky130_fd_sc_hs__fill_8 FILLER_137_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_137_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_137_423 ();
 sky130_fd_sc_hs__fill_1 FILLER_137_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_137_438 ();
 sky130_fd_sc_hs__fill_4 FILLER_137_446 ();
 sky130_fd_sc_hs__fill_2 FILLER_137_450 ();
 sky130_fd_sc_hs__fill_8 FILLER_137_456 ();
 sky130_fd_sc_hs__fill_2 FILLER_137_465 ();
 sky130_fd_sc_hs__fill_4 FILLER_137_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_137_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_137_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_137_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_138_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_138_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_138_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_138_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_138_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_138_38 ();
 sky130_fd_sc_hs__fill_4 FILLER_138_46 ();
 sky130_fd_sc_hs__fill_2 FILLER_138_50 ();
 sky130_fd_sc_hs__fill_4 FILLER_138_73 ();
 sky130_fd_sc_hs__fill_2 FILLER_138_77 ();
 sky130_fd_sc_hs__fill_1 FILLER_138_82 ();
 sky130_fd_sc_hs__fill_1 FILLER_138_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_138_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_138_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_138_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_138_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_138_120 ();
 sky130_fd_sc_hs__fill_2 FILLER_138_128 ();
 sky130_fd_sc_hs__fill_1 FILLER_138_130 ();
 sky130_fd_sc_hs__fill_2 FILLER_138_135 ();
 sky130_fd_sc_hs__fill_1 FILLER_138_137 ();
 sky130_fd_sc_hs__fill_8 FILLER_138_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_138_154 ();
 sky130_fd_sc_hs__fill_1 FILLER_138_162 ();
 sky130_fd_sc_hs__fill_4 FILLER_138_198 ();
 sky130_fd_sc_hs__fill_1 FILLER_138_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_138_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_138_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_138_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_138_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_138_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_138_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_138_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_138_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_138_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_138_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_138_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_138_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_138_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_138_302 ();
 sky130_fd_sc_hs__fill_8 FILLER_138_310 ();
 sky130_fd_sc_hs__fill_1 FILLER_138_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_138_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_138_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_138_350 ();
 sky130_fd_sc_hs__fill_8 FILLER_138_358 ();
 sky130_fd_sc_hs__fill_8 FILLER_138_366 ();
 sky130_fd_sc_hs__fill_2 FILLER_138_374 ();
 sky130_fd_sc_hs__fill_1 FILLER_138_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_138_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_138_386 ();
 sky130_fd_sc_hs__fill_4 FILLER_138_394 ();
 sky130_fd_sc_hs__fill_2 FILLER_138_398 ();
 sky130_fd_sc_hs__fill_1 FILLER_138_400 ();
 sky130_fd_sc_hs__fill_8 FILLER_138_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_138_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_138_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_138_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_138_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_138_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_138_452 ();
 sky130_fd_sc_hs__fill_4 FILLER_138_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_138_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_138_481 ();
 sky130_fd_sc_hs__fill_4 FILLER_138_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_138_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_138_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_138_510 ();
 sky130_fd_sc_hs__fill_4 FILLER_138_518 ();
 sky130_fd_sc_hs__fill_2 FILLER_138_522 ();
 sky130_fd_sc_hs__fill_8 FILLER_139_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_139_8 ();
 sky130_fd_sc_hs__fill_4 FILLER_139_16 ();
 sky130_fd_sc_hs__fill_2 FILLER_139_20 ();
 sky130_fd_sc_hs__fill_1 FILLER_139_22 ();
 sky130_fd_sc_hs__fill_8 FILLER_139_43 ();
 sky130_fd_sc_hs__fill_4 FILLER_139_51 ();
 sky130_fd_sc_hs__fill_2 FILLER_139_55 ();
 sky130_fd_sc_hs__fill_1 FILLER_139_57 ();
 sky130_fd_sc_hs__fill_2 FILLER_139_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_139_69 ();
 sky130_fd_sc_hs__fill_8 FILLER_139_77 ();
 sky130_fd_sc_hs__fill_8 FILLER_139_85 ();
 sky130_fd_sc_hs__fill_8 FILLER_139_93 ();
 sky130_fd_sc_hs__fill_8 FILLER_139_101 ();
 sky130_fd_sc_hs__fill_4 FILLER_139_109 ();
 sky130_fd_sc_hs__fill_2 FILLER_139_113 ();
 sky130_fd_sc_hs__fill_1 FILLER_139_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_139_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_139_125 ();
 sky130_fd_sc_hs__fill_4 FILLER_139_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_139_140 ();
 sky130_fd_sc_hs__fill_8 FILLER_139_148 ();
 sky130_fd_sc_hs__fill_8 FILLER_139_156 ();
 sky130_fd_sc_hs__fill_8 FILLER_139_164 ();
 sky130_fd_sc_hs__fill_2 FILLER_139_172 ();
 sky130_fd_sc_hs__fill_8 FILLER_139_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_139_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_139_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_139_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_139_207 ();
 sky130_fd_sc_hs__fill_4 FILLER_139_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_139_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_139_241 ();
 sky130_fd_sc_hs__fill_1 FILLER_139_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_139_263 ();
 sky130_fd_sc_hs__fill_8 FILLER_139_271 ();
 sky130_fd_sc_hs__fill_8 FILLER_139_279 ();
 sky130_fd_sc_hs__fill_2 FILLER_139_287 ();
 sky130_fd_sc_hs__fill_1 FILLER_139_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_139_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_139_299 ();
 sky130_fd_sc_hs__fill_4 FILLER_139_307 ();
 sky130_fd_sc_hs__fill_2 FILLER_139_311 ();
 sky130_fd_sc_hs__fill_1 FILLER_139_313 ();
 sky130_fd_sc_hs__fill_8 FILLER_139_323 ();
 sky130_fd_sc_hs__fill_1 FILLER_139_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_139_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_139_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_139_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_139_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_139_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_139_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_139_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_139_405 ();
 sky130_fd_sc_hs__fill_1 FILLER_139_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_139_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_139_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_139_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_139_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_139_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_139_481 ();
 sky130_fd_sc_hs__fill_1 FILLER_139_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_139_498 ();
 sky130_fd_sc_hs__fill_8 FILLER_139_506 ();
 sky130_fd_sc_hs__fill_2 FILLER_139_514 ();
 sky130_fd_sc_hs__fill_2 FILLER_139_519 ();
 sky130_fd_sc_hs__fill_1 FILLER_139_521 ();
 sky130_fd_sc_hs__fill_1 FILLER_139_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_139_532 ();
 sky130_fd_sc_hs__fill_8 FILLER_140_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_140_8 ();
 sky130_fd_sc_hs__fill_4 FILLER_140_16 ();
 sky130_fd_sc_hs__fill_1 FILLER_140_20 ();
 sky130_fd_sc_hs__fill_4 FILLER_140_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_140_49 ();
 sky130_fd_sc_hs__fill_8 FILLER_140_57 ();
 sky130_fd_sc_hs__fill_8 FILLER_140_65 ();
 sky130_fd_sc_hs__fill_8 FILLER_140_73 ();
 sky130_fd_sc_hs__fill_4 FILLER_140_81 ();
 sky130_fd_sc_hs__fill_2 FILLER_140_85 ();
 sky130_fd_sc_hs__fill_8 FILLER_140_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_140_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_140_108 ();
 sky130_fd_sc_hs__fill_8 FILLER_140_116 ();
 sky130_fd_sc_hs__fill_4 FILLER_140_124 ();
 sky130_fd_sc_hs__fill_1 FILLER_140_128 ();
 sky130_fd_sc_hs__fill_4 FILLER_140_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_140_146 ();
 sky130_fd_sc_hs__fill_4 FILLER_140_154 ();
 sky130_fd_sc_hs__fill_2 FILLER_140_158 ();
 sky130_fd_sc_hs__fill_4 FILLER_140_196 ();
 sky130_fd_sc_hs__fill_2 FILLER_140_200 ();
 sky130_fd_sc_hs__fill_1 FILLER_140_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_140_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_140_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_140_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_140_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_140_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_140_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_140_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_140_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_140_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_140_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_140_286 ();
 sky130_fd_sc_hs__fill_4 FILLER_140_294 ();
 sky130_fd_sc_hs__fill_1 FILLER_140_298 ();
 sky130_fd_sc_hs__fill_8 FILLER_140_310 ();
 sky130_fd_sc_hs__fill_1 FILLER_140_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_140_341 ();
 sky130_fd_sc_hs__fill_8 FILLER_140_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_140_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_140_365 ();
 sky130_fd_sc_hs__fill_4 FILLER_140_373 ();
 sky130_fd_sc_hs__fill_2 FILLER_140_378 ();
 sky130_fd_sc_hs__fill_1 FILLER_140_398 ();
 sky130_fd_sc_hs__fill_8 FILLER_140_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_140_410 ();
 sky130_fd_sc_hs__fill_4 FILLER_140_418 ();
 sky130_fd_sc_hs__fill_2 FILLER_140_422 ();
 sky130_fd_sc_hs__fill_1 FILLER_140_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_140_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_140_444 ();
 sky130_fd_sc_hs__fill_2 FILLER_140_452 ();
 sky130_fd_sc_hs__fill_1 FILLER_140_454 ();
 sky130_fd_sc_hs__fill_8 FILLER_140_467 ();
 sky130_fd_sc_hs__fill_8 FILLER_140_475 ();
 sky130_fd_sc_hs__fill_8 FILLER_140_483 ();
 sky130_fd_sc_hs__fill_2 FILLER_140_491 ();
 sky130_fd_sc_hs__fill_8 FILLER_140_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_140_502 ();
 sky130_fd_sc_hs__fill_1 FILLER_140_510 ();
 sky130_fd_sc_hs__fill_4 FILLER_140_521 ();
 sky130_fd_sc_hs__fill_1 FILLER_140_525 ();
 sky130_fd_sc_hs__fill_2 FILLER_140_537 ();
 sky130_fd_sc_hs__fill_1 FILLER_140_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_141_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_141_8 ();
 sky130_fd_sc_hs__fill_2 FILLER_141_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_141_26 ();
 sky130_fd_sc_hs__fill_2 FILLER_141_34 ();
 sky130_fd_sc_hs__fill_1 FILLER_141_36 ();
 sky130_fd_sc_hs__fill_8 FILLER_141_50 ();
 sky130_fd_sc_hs__fill_8 FILLER_141_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_141_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_141_75 ();
 sky130_fd_sc_hs__fill_2 FILLER_141_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_141_106 ();
 sky130_fd_sc_hs__fill_2 FILLER_141_114 ();
 sky130_fd_sc_hs__fill_8 FILLER_141_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_141_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_141_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_141_162 ();
 sky130_fd_sc_hs__fill_4 FILLER_141_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_141_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_141_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_141_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_141_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_141_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_141_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_141_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_141_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_141_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_141_241 ();
 sky130_fd_sc_hs__fill_2 FILLER_141_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_141_269 ();
 sky130_fd_sc_hs__fill_8 FILLER_141_277 ();
 sky130_fd_sc_hs__fill_4 FILLER_141_285 ();
 sky130_fd_sc_hs__fill_1 FILLER_141_289 ();
 sky130_fd_sc_hs__fill_2 FILLER_141_291 ();
 sky130_fd_sc_hs__fill_1 FILLER_141_293 ();
 sky130_fd_sc_hs__fill_4 FILLER_141_311 ();
 sky130_fd_sc_hs__fill_2 FILLER_141_315 ();
 sky130_fd_sc_hs__fill_1 FILLER_141_317 ();
 sky130_fd_sc_hs__fill_8 FILLER_141_335 ();
 sky130_fd_sc_hs__fill_4 FILLER_141_343 ();
 sky130_fd_sc_hs__fill_1 FILLER_141_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_141_349 ();
 sky130_fd_sc_hs__fill_4 FILLER_141_357 ();
 sky130_fd_sc_hs__fill_1 FILLER_141_361 ();
 sky130_fd_sc_hs__fill_1 FILLER_141_369 ();
 sky130_fd_sc_hs__fill_8 FILLER_141_380 ();
 sky130_fd_sc_hs__fill_2 FILLER_141_388 ();
 sky130_fd_sc_hs__fill_8 FILLER_141_395 ();
 sky130_fd_sc_hs__fill_2 FILLER_141_403 ();
 sky130_fd_sc_hs__fill_1 FILLER_141_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_141_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_141_415 ();
 sky130_fd_sc_hs__fill_1 FILLER_141_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_141_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_141_442 ();
 sky130_fd_sc_hs__fill_2 FILLER_141_450 ();
 sky130_fd_sc_hs__fill_2 FILLER_141_461 ();
 sky130_fd_sc_hs__fill_1 FILLER_141_463 ();
 sky130_fd_sc_hs__fill_4 FILLER_141_488 ();
 sky130_fd_sc_hs__fill_2 FILLER_141_492 ();
 sky130_fd_sc_hs__fill_4 FILLER_141_502 ();
 sky130_fd_sc_hs__fill_1 FILLER_141_506 ();
 sky130_fd_sc_hs__fill_4 FILLER_141_517 ();
 sky130_fd_sc_hs__fill_1 FILLER_141_521 ();
 sky130_fd_sc_hs__fill_4 FILLER_141_533 ();
 sky130_fd_sc_hs__fill_2 FILLER_141_537 ();
 sky130_fd_sc_hs__fill_1 FILLER_141_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_142_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_142_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_142_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_142_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_142_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_142_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_142_52 ();
 sky130_fd_sc_hs__fill_8 FILLER_142_60 ();
 sky130_fd_sc_hs__fill_8 FILLER_142_68 ();
 sky130_fd_sc_hs__fill_8 FILLER_142_76 ();
 sky130_fd_sc_hs__fill_2 FILLER_142_84 ();
 sky130_fd_sc_hs__fill_1 FILLER_142_86 ();
 sky130_fd_sc_hs__fill_1 FILLER_142_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_142_94 ();
 sky130_fd_sc_hs__fill_8 FILLER_142_102 ();
 sky130_fd_sc_hs__fill_4 FILLER_142_110 ();
 sky130_fd_sc_hs__fill_2 FILLER_142_114 ();
 sky130_fd_sc_hs__fill_2 FILLER_142_128 ();
 sky130_fd_sc_hs__fill_1 FILLER_142_130 ();
 sky130_fd_sc_hs__fill_4 FILLER_142_135 ();
 sky130_fd_sc_hs__fill_1 FILLER_142_139 ();
 sky130_fd_sc_hs__fill_1 FILLER_142_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_142_153 ();
 sky130_fd_sc_hs__fill_8 FILLER_142_161 ();
 sky130_fd_sc_hs__fill_8 FILLER_142_169 ();
 sky130_fd_sc_hs__fill_8 FILLER_142_177 ();
 sky130_fd_sc_hs__fill_8 FILLER_142_185 ();
 sky130_fd_sc_hs__fill_8 FILLER_142_193 ();
 sky130_fd_sc_hs__fill_2 FILLER_142_201 ();
 sky130_fd_sc_hs__fill_4 FILLER_142_204 ();
 sky130_fd_sc_hs__fill_1 FILLER_142_208 ();
 sky130_fd_sc_hs__fill_2 FILLER_142_239 ();
 sky130_fd_sc_hs__fill_1 FILLER_142_241 ();
 sky130_fd_sc_hs__fill_2 FILLER_142_262 ();
 sky130_fd_sc_hs__fill_2 FILLER_142_272 ();
 sky130_fd_sc_hs__fill_4 FILLER_142_306 ();
 sky130_fd_sc_hs__fill_8 FILLER_142_320 ();
 sky130_fd_sc_hs__fill_2 FILLER_142_328 ();
 sky130_fd_sc_hs__fill_1 FILLER_142_330 ();
 sky130_fd_sc_hs__fill_8 FILLER_142_340 ();
 sky130_fd_sc_hs__fill_8 FILLER_142_348 ();
 sky130_fd_sc_hs__fill_8 FILLER_142_356 ();
 sky130_fd_sc_hs__fill_8 FILLER_142_364 ();
 sky130_fd_sc_hs__fill_4 FILLER_142_372 ();
 sky130_fd_sc_hs__fill_1 FILLER_142_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_142_378 ();
 sky130_fd_sc_hs__fill_4 FILLER_142_386 ();
 sky130_fd_sc_hs__fill_2 FILLER_142_400 ();
 sky130_fd_sc_hs__fill_1 FILLER_142_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_142_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_142_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_142_478 ();
 sky130_fd_sc_hs__fill_4 FILLER_142_486 ();
 sky130_fd_sc_hs__fill_2 FILLER_142_490 ();
 sky130_fd_sc_hs__fill_1 FILLER_142_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_142_494 ();
 sky130_fd_sc_hs__fill_2 FILLER_142_502 ();
 sky130_fd_sc_hs__fill_1 FILLER_142_504 ();
 sky130_fd_sc_hs__fill_4 FILLER_142_535 ();
 sky130_fd_sc_hs__fill_1 FILLER_142_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_143_0 ();
 sky130_fd_sc_hs__fill_2 FILLER_143_8 ();
 sky130_fd_sc_hs__fill_1 FILLER_143_10 ();
 sky130_fd_sc_hs__fill_8 FILLER_143_19 ();
 sky130_fd_sc_hs__fill_8 FILLER_143_27 ();
 sky130_fd_sc_hs__fill_8 FILLER_143_35 ();
 sky130_fd_sc_hs__fill_8 FILLER_143_43 ();
 sky130_fd_sc_hs__fill_4 FILLER_143_51 ();
 sky130_fd_sc_hs__fill_2 FILLER_143_55 ();
 sky130_fd_sc_hs__fill_1 FILLER_143_57 ();
 sky130_fd_sc_hs__fill_8 FILLER_143_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_143_67 ();
 sky130_fd_sc_hs__fill_2 FILLER_143_75 ();
 sky130_fd_sc_hs__fill_1 FILLER_143_77 ();
 sky130_fd_sc_hs__fill_4 FILLER_143_101 ();
 sky130_fd_sc_hs__fill_4 FILLER_143_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_143_163 ();
 sky130_fd_sc_hs__fill_2 FILLER_143_171 ();
 sky130_fd_sc_hs__fill_1 FILLER_143_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_143_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_143_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_143_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_143_199 ();
 sky130_fd_sc_hs__fill_2 FILLER_143_207 ();
 sky130_fd_sc_hs__fill_4 FILLER_143_226 ();
 sky130_fd_sc_hs__fill_2 FILLER_143_230 ();
 sky130_fd_sc_hs__fill_8 FILLER_143_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_143_241 ();
 sky130_fd_sc_hs__fill_4 FILLER_143_249 ();
 sky130_fd_sc_hs__fill_4 FILLER_143_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_143_278 ();
 sky130_fd_sc_hs__fill_4 FILLER_143_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_143_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_143_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_143_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_143_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_143_323 ();
 sky130_fd_sc_hs__fill_2 FILLER_143_331 ();
 sky130_fd_sc_hs__fill_4 FILLER_143_343 ();
 sky130_fd_sc_hs__fill_1 FILLER_143_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_143_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_143_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_143_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_143_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_143_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_143_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_143_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_143_405 ();
 sky130_fd_sc_hs__fill_4 FILLER_143_407 ();
 sky130_fd_sc_hs__fill_2 FILLER_143_411 ();
 sky130_fd_sc_hs__fill_1 FILLER_143_413 ();
 sky130_fd_sc_hs__fill_8 FILLER_143_421 ();
 sky130_fd_sc_hs__fill_8 FILLER_143_429 ();
 sky130_fd_sc_hs__fill_8 FILLER_143_437 ();
 sky130_fd_sc_hs__fill_8 FILLER_143_445 ();
 sky130_fd_sc_hs__fill_1 FILLER_143_453 ();
 sky130_fd_sc_hs__fill_4 FILLER_143_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_143_477 ();
 sky130_fd_sc_hs__fill_8 FILLER_143_485 ();
 sky130_fd_sc_hs__fill_4 FILLER_143_493 ();
 sky130_fd_sc_hs__fill_1 FILLER_143_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_143_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_143_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_144_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_144_8 ();
 sky130_fd_sc_hs__fill_4 FILLER_144_16 ();
 sky130_fd_sc_hs__fill_1 FILLER_144_20 ();
 sky130_fd_sc_hs__fill_8 FILLER_144_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_144_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_144_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_144_54 ();
 sky130_fd_sc_hs__fill_2 FILLER_144_62 ();
 sky130_fd_sc_hs__fill_1 FILLER_144_64 ();
 sky130_fd_sc_hs__fill_4 FILLER_144_77 ();
 sky130_fd_sc_hs__fill_2 FILLER_144_81 ();
 sky130_fd_sc_hs__fill_8 FILLER_144_100 ();
 sky130_fd_sc_hs__fill_8 FILLER_144_108 ();
 sky130_fd_sc_hs__fill_8 FILLER_144_116 ();
 sky130_fd_sc_hs__fill_8 FILLER_144_124 ();
 sky130_fd_sc_hs__fill_8 FILLER_144_132 ();
 sky130_fd_sc_hs__fill_4 FILLER_144_140 ();
 sky130_fd_sc_hs__fill_1 FILLER_144_144 ();
 sky130_fd_sc_hs__fill_1 FILLER_144_146 ();
 sky130_fd_sc_hs__fill_1 FILLER_144_160 ();
 sky130_fd_sc_hs__fill_2 FILLER_144_187 ();
 sky130_fd_sc_hs__fill_1 FILLER_144_189 ();
 sky130_fd_sc_hs__fill_8 FILLER_144_193 ();
 sky130_fd_sc_hs__fill_2 FILLER_144_201 ();
 sky130_fd_sc_hs__fill_2 FILLER_144_209 ();
 sky130_fd_sc_hs__fill_8 FILLER_144_228 ();
 sky130_fd_sc_hs__fill_1 FILLER_144_236 ();
 sky130_fd_sc_hs__fill_4 FILLER_144_256 ();
 sky130_fd_sc_hs__fill_1 FILLER_144_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_144_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_144_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_144_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_144_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_144_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_144_302 ();
 sky130_fd_sc_hs__fill_8 FILLER_144_310 ();
 sky130_fd_sc_hs__fill_1 FILLER_144_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_144_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_144_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_144_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_144_344 ();
 sky130_fd_sc_hs__fill_2 FILLER_144_352 ();
 sky130_fd_sc_hs__fill_1 FILLER_144_354 ();
 sky130_fd_sc_hs__fill_8 FILLER_144_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_144_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_144_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_144_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_144_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_144_418 ();
 sky130_fd_sc_hs__fill_2 FILLER_144_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_144_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_144_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_144_444 ();
 sky130_fd_sc_hs__fill_2 FILLER_144_491 ();
 sky130_fd_sc_hs__fill_4 FILLER_144_494 ();
 sky130_fd_sc_hs__fill_2 FILLER_144_498 ();
 sky130_fd_sc_hs__fill_1 FILLER_144_500 ();
 sky130_fd_sc_hs__fill_2 FILLER_144_509 ();
 sky130_fd_sc_hs__fill_8 FILLER_144_523 ();
 sky130_fd_sc_hs__fill_1 FILLER_144_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_145_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_145_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_145_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_145_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_145_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_145_45 ();
 sky130_fd_sc_hs__fill_4 FILLER_145_53 ();
 sky130_fd_sc_hs__fill_1 FILLER_145_57 ();
 sky130_fd_sc_hs__fill_8 FILLER_145_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_145_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_145_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_145_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_145_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_145_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_145_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_145_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_145_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_145_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_145_133 ();
 sky130_fd_sc_hs__fill_4 FILLER_145_141 ();
 sky130_fd_sc_hs__fill_1 FILLER_145_145 ();
 sky130_fd_sc_hs__fill_1 FILLER_145_152 ();
 sky130_fd_sc_hs__fill_1 FILLER_145_157 ();
 sky130_fd_sc_hs__fill_4 FILLER_145_168 ();
 sky130_fd_sc_hs__fill_2 FILLER_145_172 ();
 sky130_fd_sc_hs__fill_2 FILLER_145_175 ();
 sky130_fd_sc_hs__fill_2 FILLER_145_207 ();
 sky130_fd_sc_hs__fill_2 FILLER_145_225 ();
 sky130_fd_sc_hs__fill_1 FILLER_145_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_145_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_145_252 ();
 sky130_fd_sc_hs__fill_4 FILLER_145_260 ();
 sky130_fd_sc_hs__fill_2 FILLER_145_264 ();
 sky130_fd_sc_hs__fill_1 FILLER_145_266 ();
 sky130_fd_sc_hs__fill_8 FILLER_145_279 ();
 sky130_fd_sc_hs__fill_2 FILLER_145_287 ();
 sky130_fd_sc_hs__fill_1 FILLER_145_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_145_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_145_299 ();
 sky130_fd_sc_hs__fill_4 FILLER_145_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_145_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_145_336 ();
 sky130_fd_sc_hs__fill_4 FILLER_145_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_145_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_145_357 ();
 sky130_fd_sc_hs__fill_4 FILLER_145_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_145_387 ();
 sky130_fd_sc_hs__fill_8 FILLER_145_395 ();
 sky130_fd_sc_hs__fill_2 FILLER_145_403 ();
 sky130_fd_sc_hs__fill_1 FILLER_145_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_145_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_145_415 ();
 sky130_fd_sc_hs__fill_4 FILLER_145_423 ();
 sky130_fd_sc_hs__fill_1 FILLER_145_427 ();
 sky130_fd_sc_hs__fill_8 FILLER_145_432 ();
 sky130_fd_sc_hs__fill_8 FILLER_145_440 ();
 sky130_fd_sc_hs__fill_8 FILLER_145_452 ();
 sky130_fd_sc_hs__fill_4 FILLER_145_460 ();
 sky130_fd_sc_hs__fill_1 FILLER_145_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_145_479 ();
 sky130_fd_sc_hs__fill_8 FILLER_145_487 ();
 sky130_fd_sc_hs__fill_8 FILLER_145_495 ();
 sky130_fd_sc_hs__fill_2 FILLER_145_503 ();
 sky130_fd_sc_hs__fill_4 FILLER_145_517 ();
 sky130_fd_sc_hs__fill_1 FILLER_145_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_145_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_145_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_145_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_146_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_146_8 ();
 sky130_fd_sc_hs__fill_4 FILLER_146_16 ();
 sky130_fd_sc_hs__fill_1 FILLER_146_20 ();
 sky130_fd_sc_hs__fill_8 FILLER_146_30 ();
 sky130_fd_sc_hs__fill_2 FILLER_146_38 ();
 sky130_fd_sc_hs__fill_1 FILLER_146_40 ();
 sky130_fd_sc_hs__fill_4 FILLER_146_81 ();
 sky130_fd_sc_hs__fill_2 FILLER_146_85 ();
 sky130_fd_sc_hs__fill_8 FILLER_146_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_146_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_146_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_146_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_146_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_146_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_146_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_146_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_146_146 ();
 sky130_fd_sc_hs__fill_2 FILLER_146_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_146_162 ();
 sky130_fd_sc_hs__fill_2 FILLER_146_170 ();
 sky130_fd_sc_hs__fill_1 FILLER_146_172 ();
 sky130_fd_sc_hs__fill_4 FILLER_146_199 ();
 sky130_fd_sc_hs__fill_1 FILLER_146_216 ();
 sky130_fd_sc_hs__fill_4 FILLER_146_224 ();
 sky130_fd_sc_hs__fill_1 FILLER_146_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_146_247 ();
 sky130_fd_sc_hs__fill_4 FILLER_146_255 ();
 sky130_fd_sc_hs__fill_2 FILLER_146_259 ();
 sky130_fd_sc_hs__fill_8 FILLER_146_262 ();
 sky130_fd_sc_hs__fill_4 FILLER_146_270 ();
 sky130_fd_sc_hs__fill_1 FILLER_146_274 ();
 sky130_fd_sc_hs__fill_8 FILLER_146_287 ();
 sky130_fd_sc_hs__fill_8 FILLER_146_295 ();
 sky130_fd_sc_hs__fill_8 FILLER_146_303 ();
 sky130_fd_sc_hs__fill_4 FILLER_146_311 ();
 sky130_fd_sc_hs__fill_1 FILLER_146_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_146_320 ();
 sky130_fd_sc_hs__fill_4 FILLER_146_336 ();
 sky130_fd_sc_hs__fill_2 FILLER_146_340 ();
 sky130_fd_sc_hs__fill_1 FILLER_146_342 ();
 sky130_fd_sc_hs__fill_8 FILLER_146_364 ();
 sky130_fd_sc_hs__fill_4 FILLER_146_372 ();
 sky130_fd_sc_hs__fill_1 FILLER_146_376 ();
 sky130_fd_sc_hs__fill_2 FILLER_146_378 ();
 sky130_fd_sc_hs__fill_1 FILLER_146_380 ();
 sky130_fd_sc_hs__fill_1 FILLER_146_390 ();
 sky130_fd_sc_hs__fill_2 FILLER_146_416 ();
 sky130_fd_sc_hs__fill_1 FILLER_146_418 ();
 sky130_fd_sc_hs__fill_2 FILLER_146_436 ();
 sky130_fd_sc_hs__fill_1 FILLER_146_438 ();
 sky130_fd_sc_hs__fill_2 FILLER_146_460 ();
 sky130_fd_sc_hs__fill_1 FILLER_146_462 ();
 sky130_fd_sc_hs__fill_8 FILLER_146_467 ();
 sky130_fd_sc_hs__fill_2 FILLER_146_475 ();
 sky130_fd_sc_hs__fill_1 FILLER_146_477 ();
 sky130_fd_sc_hs__fill_4 FILLER_146_487 ();
 sky130_fd_sc_hs__fill_2 FILLER_146_491 ();
 sky130_fd_sc_hs__fill_8 FILLER_146_517 ();
 sky130_fd_sc_hs__fill_2 FILLER_146_525 ();
 sky130_fd_sc_hs__fill_1 FILLER_146_527 ();
 sky130_fd_sc_hs__fill_4 FILLER_146_536 ();
 sky130_fd_sc_hs__fill_8 FILLER_147_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_147_8 ();
 sky130_fd_sc_hs__fill_4 FILLER_147_16 ();
 sky130_fd_sc_hs__fill_2 FILLER_147_20 ();
 sky130_fd_sc_hs__fill_4 FILLER_147_40 ();
 sky130_fd_sc_hs__fill_1 FILLER_147_44 ();
 sky130_fd_sc_hs__fill_8 FILLER_147_59 ();
 sky130_fd_sc_hs__fill_2 FILLER_147_67 ();
 sky130_fd_sc_hs__fill_2 FILLER_147_90 ();
 sky130_fd_sc_hs__fill_2 FILLER_147_113 ();
 sky130_fd_sc_hs__fill_1 FILLER_147_115 ();
 sky130_fd_sc_hs__fill_2 FILLER_147_117 ();
 sky130_fd_sc_hs__fill_2 FILLER_147_137 ();
 sky130_fd_sc_hs__fill_1 FILLER_147_139 ();
 sky130_fd_sc_hs__fill_2 FILLER_147_156 ();
 sky130_fd_sc_hs__fill_1 FILLER_147_158 ();
 sky130_fd_sc_hs__fill_1 FILLER_147_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_147_175 ();
 sky130_fd_sc_hs__fill_4 FILLER_147_183 ();
 sky130_fd_sc_hs__fill_2 FILLER_147_187 ();
 sky130_fd_sc_hs__fill_8 FILLER_147_200 ();
 sky130_fd_sc_hs__fill_8 FILLER_147_208 ();
 sky130_fd_sc_hs__fill_4 FILLER_147_216 ();
 sky130_fd_sc_hs__fill_2 FILLER_147_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_147_251 ();
 sky130_fd_sc_hs__fill_8 FILLER_147_259 ();
 sky130_fd_sc_hs__fill_8 FILLER_147_267 ();
 sky130_fd_sc_hs__fill_8 FILLER_147_275 ();
 sky130_fd_sc_hs__fill_4 FILLER_147_283 ();
 sky130_fd_sc_hs__fill_2 FILLER_147_287 ();
 sky130_fd_sc_hs__fill_1 FILLER_147_289 ();
 sky130_fd_sc_hs__fill_4 FILLER_147_291 ();
 sky130_fd_sc_hs__fill_2 FILLER_147_295 ();
 sky130_fd_sc_hs__fill_1 FILLER_147_297 ();
 sky130_fd_sc_hs__fill_8 FILLER_147_314 ();
 sky130_fd_sc_hs__fill_4 FILLER_147_322 ();
 sky130_fd_sc_hs__fill_1 FILLER_147_326 ();
 sky130_fd_sc_hs__fill_4 FILLER_147_343 ();
 sky130_fd_sc_hs__fill_1 FILLER_147_347 ();
 sky130_fd_sc_hs__fill_2 FILLER_147_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_147_395 ();
 sky130_fd_sc_hs__fill_2 FILLER_147_403 ();
 sky130_fd_sc_hs__fill_1 FILLER_147_405 ();
 sky130_fd_sc_hs__fill_4 FILLER_147_407 ();
 sky130_fd_sc_hs__fill_1 FILLER_147_411 ();
 sky130_fd_sc_hs__fill_4 FILLER_147_428 ();
 sky130_fd_sc_hs__fill_2 FILLER_147_450 ();
 sky130_fd_sc_hs__fill_1 FILLER_147_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_147_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_147_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_147_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_147_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_147_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_147_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_147_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_148_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_148_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_148_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_148_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_148_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_148_38 ();
 sky130_fd_sc_hs__fill_4 FILLER_148_46 ();
 sky130_fd_sc_hs__fill_2 FILLER_148_50 ();
 sky130_fd_sc_hs__fill_1 FILLER_148_52 ();
 sky130_fd_sc_hs__fill_1 FILLER_148_65 ();
 sky130_fd_sc_hs__fill_4 FILLER_148_88 ();
 sky130_fd_sc_hs__fill_2 FILLER_148_92 ();
 sky130_fd_sc_hs__fill_8 FILLER_148_102 ();
 sky130_fd_sc_hs__fill_8 FILLER_148_110 ();
 sky130_fd_sc_hs__fill_4 FILLER_148_118 ();
 sky130_fd_sc_hs__fill_1 FILLER_148_122 ();
 sky130_fd_sc_hs__fill_2 FILLER_148_143 ();
 sky130_fd_sc_hs__fill_2 FILLER_148_146 ();
 sky130_fd_sc_hs__fill_4 FILLER_148_152 ();
 sky130_fd_sc_hs__fill_2 FILLER_148_156 ();
 sky130_fd_sc_hs__fill_1 FILLER_148_158 ();
 sky130_fd_sc_hs__fill_8 FILLER_148_164 ();
 sky130_fd_sc_hs__fill_8 FILLER_148_172 ();
 sky130_fd_sc_hs__fill_8 FILLER_148_180 ();
 sky130_fd_sc_hs__fill_8 FILLER_148_188 ();
 sky130_fd_sc_hs__fill_4 FILLER_148_196 ();
 sky130_fd_sc_hs__fill_2 FILLER_148_200 ();
 sky130_fd_sc_hs__fill_1 FILLER_148_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_148_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_148_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_148_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_148_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_148_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_148_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_148_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_148_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_148_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_148_270 ();
 sky130_fd_sc_hs__fill_1 FILLER_148_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_148_296 ();
 sky130_fd_sc_hs__fill_8 FILLER_148_304 ();
 sky130_fd_sc_hs__fill_4 FILLER_148_312 ();
 sky130_fd_sc_hs__fill_2 FILLER_148_316 ();
 sky130_fd_sc_hs__fill_1 FILLER_148_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_148_332 ();
 sky130_fd_sc_hs__fill_4 FILLER_148_340 ();
 sky130_fd_sc_hs__fill_2 FILLER_148_344 ();
 sky130_fd_sc_hs__fill_1 FILLER_148_346 ();
 sky130_fd_sc_hs__fill_4 FILLER_148_370 ();
 sky130_fd_sc_hs__fill_2 FILLER_148_374 ();
 sky130_fd_sc_hs__fill_1 FILLER_148_376 ();
 sky130_fd_sc_hs__fill_4 FILLER_148_378 ();
 sky130_fd_sc_hs__fill_1 FILLER_148_382 ();
 sky130_fd_sc_hs__fill_8 FILLER_148_413 ();
 sky130_fd_sc_hs__fill_8 FILLER_148_421 ();
 sky130_fd_sc_hs__fill_4 FILLER_148_429 ();
 sky130_fd_sc_hs__fill_2 FILLER_148_433 ();
 sky130_fd_sc_hs__fill_4 FILLER_148_436 ();
 sky130_fd_sc_hs__fill_2 FILLER_148_443 ();
 sky130_fd_sc_hs__fill_8 FILLER_148_451 ();
 sky130_fd_sc_hs__fill_8 FILLER_148_459 ();
 sky130_fd_sc_hs__fill_8 FILLER_148_467 ();
 sky130_fd_sc_hs__fill_8 FILLER_148_475 ();
 sky130_fd_sc_hs__fill_8 FILLER_148_483 ();
 sky130_fd_sc_hs__fill_2 FILLER_148_491 ();
 sky130_fd_sc_hs__fill_8 FILLER_148_501 ();
 sky130_fd_sc_hs__fill_4 FILLER_148_509 ();
 sky130_fd_sc_hs__fill_2 FILLER_148_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_148_515 ();
 sky130_fd_sc_hs__fill_4 FILLER_148_524 ();
 sky130_fd_sc_hs__fill_1 FILLER_148_528 ();
 sky130_fd_sc_hs__fill_2 FILLER_148_537 ();
 sky130_fd_sc_hs__fill_1 FILLER_148_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_149_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_149_8 ();
 sky130_fd_sc_hs__fill_1 FILLER_149_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_149_47 ();
 sky130_fd_sc_hs__fill_2 FILLER_149_55 ();
 sky130_fd_sc_hs__fill_1 FILLER_149_57 ();
 sky130_fd_sc_hs__fill_8 FILLER_149_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_149_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_149_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_149_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_149_91 ();
 sky130_fd_sc_hs__fill_4 FILLER_149_99 ();
 sky130_fd_sc_hs__fill_2 FILLER_149_103 ();
 sky130_fd_sc_hs__fill_8 FILLER_149_117 ();
 sky130_fd_sc_hs__fill_2 FILLER_149_128 ();
 sky130_fd_sc_hs__fill_2 FILLER_149_134 ();
 sky130_fd_sc_hs__fill_2 FILLER_149_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_149_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_149_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_149_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_149_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_149_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_149_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_149_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_149_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_149_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_149_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_149_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_149_257 ();
 sky130_fd_sc_hs__fill_2 FILLER_149_265 ();
 sky130_fd_sc_hs__fill_1 FILLER_149_267 ();
 sky130_fd_sc_hs__fill_8 FILLER_149_276 ();
 sky130_fd_sc_hs__fill_4 FILLER_149_284 ();
 sky130_fd_sc_hs__fill_2 FILLER_149_288 ();
 sky130_fd_sc_hs__fill_1 FILLER_149_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_149_309 ();
 sky130_fd_sc_hs__fill_8 FILLER_149_317 ();
 sky130_fd_sc_hs__fill_8 FILLER_149_325 ();
 sky130_fd_sc_hs__fill_8 FILLER_149_333 ();
 sky130_fd_sc_hs__fill_4 FILLER_149_341 ();
 sky130_fd_sc_hs__fill_2 FILLER_149_345 ();
 sky130_fd_sc_hs__fill_1 FILLER_149_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_149_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_149_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_149_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_149_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_149_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_149_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_149_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_149_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_149_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_149_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_149_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_149_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_149_439 ();
 sky130_fd_sc_hs__fill_4 FILLER_149_447 ();
 sky130_fd_sc_hs__fill_1 FILLER_149_451 ();
 sky130_fd_sc_hs__fill_4 FILLER_149_465 ();
 sky130_fd_sc_hs__fill_2 FILLER_149_474 ();
 sky130_fd_sc_hs__fill_1 FILLER_149_476 ();
 sky130_fd_sc_hs__fill_4 FILLER_149_516 ();
 sky130_fd_sc_hs__fill_2 FILLER_149_520 ();
 sky130_fd_sc_hs__fill_8 FILLER_149_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_149_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_149_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_150_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_150_8 ();
 sky130_fd_sc_hs__fill_2 FILLER_150_16 ();
 sky130_fd_sc_hs__fill_2 FILLER_150_26 ();
 sky130_fd_sc_hs__fill_1 FILLER_150_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_150_35 ();
 sky130_fd_sc_hs__fill_8 FILLER_150_43 ();
 sky130_fd_sc_hs__fill_8 FILLER_150_51 ();
 sky130_fd_sc_hs__fill_8 FILLER_150_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_150_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_150_75 ();
 sky130_fd_sc_hs__fill_4 FILLER_150_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_150_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_150_96 ();
 sky130_fd_sc_hs__fill_2 FILLER_150_104 ();
 sky130_fd_sc_hs__fill_4 FILLER_150_124 ();
 sky130_fd_sc_hs__fill_2 FILLER_150_128 ();
 sky130_fd_sc_hs__fill_1 FILLER_150_130 ();
 sky130_fd_sc_hs__fill_2 FILLER_150_146 ();
 sky130_fd_sc_hs__fill_4 FILLER_150_152 ();
 sky130_fd_sc_hs__fill_2 FILLER_150_156 ();
 sky130_fd_sc_hs__fill_8 FILLER_150_163 ();
 sky130_fd_sc_hs__fill_8 FILLER_150_171 ();
 sky130_fd_sc_hs__fill_8 FILLER_150_179 ();
 sky130_fd_sc_hs__fill_8 FILLER_150_187 ();
 sky130_fd_sc_hs__fill_2 FILLER_150_200 ();
 sky130_fd_sc_hs__fill_1 FILLER_150_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_150_204 ();
 sky130_fd_sc_hs__fill_1 FILLER_150_212 ();
 sky130_fd_sc_hs__fill_4 FILLER_150_227 ();
 sky130_fd_sc_hs__fill_8 FILLER_150_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_150_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_150_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_150_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_150_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_150_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_150_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_150_302 ();
 sky130_fd_sc_hs__fill_8 FILLER_150_310 ();
 sky130_fd_sc_hs__fill_1 FILLER_150_318 ();
 sky130_fd_sc_hs__fill_4 FILLER_150_320 ();
 sky130_fd_sc_hs__fill_2 FILLER_150_324 ();
 sky130_fd_sc_hs__fill_1 FILLER_150_326 ();
 sky130_fd_sc_hs__fill_8 FILLER_150_333 ();
 sky130_fd_sc_hs__fill_8 FILLER_150_341 ();
 sky130_fd_sc_hs__fill_8 FILLER_150_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_150_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_150_365 ();
 sky130_fd_sc_hs__fill_4 FILLER_150_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_150_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_150_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_150_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_150_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_150_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_150_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_150_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_150_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_150_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_150_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_150_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_150_460 ();
 sky130_fd_sc_hs__fill_2 FILLER_150_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_150_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_150_492 ();
 sky130_fd_sc_hs__fill_1 FILLER_150_494 ();
 sky130_fd_sc_hs__fill_2 FILLER_150_538 ();
 sky130_fd_sc_hs__fill_8 FILLER_151_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_151_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_151_24 ();
 sky130_fd_sc_hs__fill_2 FILLER_151_32 ();
 sky130_fd_sc_hs__fill_1 FILLER_151_34 ();
 sky130_fd_sc_hs__fill_2 FILLER_151_55 ();
 sky130_fd_sc_hs__fill_1 FILLER_151_57 ();
 sky130_fd_sc_hs__fill_8 FILLER_151_63 ();
 sky130_fd_sc_hs__fill_8 FILLER_151_71 ();
 sky130_fd_sc_hs__fill_8 FILLER_151_79 ();
 sky130_fd_sc_hs__fill_8 FILLER_151_87 ();
 sky130_fd_sc_hs__fill_8 FILLER_151_95 ();
 sky130_fd_sc_hs__fill_8 FILLER_151_103 ();
 sky130_fd_sc_hs__fill_4 FILLER_151_111 ();
 sky130_fd_sc_hs__fill_1 FILLER_151_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_151_117 ();
 sky130_fd_sc_hs__fill_4 FILLER_151_125 ();
 sky130_fd_sc_hs__fill_1 FILLER_151_129 ();
 sky130_fd_sc_hs__fill_8 FILLER_151_142 ();
 sky130_fd_sc_hs__fill_8 FILLER_151_150 ();
 sky130_fd_sc_hs__fill_8 FILLER_151_158 ();
 sky130_fd_sc_hs__fill_8 FILLER_151_166 ();
 sky130_fd_sc_hs__fill_8 FILLER_151_175 ();
 sky130_fd_sc_hs__fill_4 FILLER_151_194 ();
 sky130_fd_sc_hs__fill_2 FILLER_151_198 ();
 sky130_fd_sc_hs__fill_1 FILLER_151_200 ();
 sky130_fd_sc_hs__fill_2 FILLER_151_216 ();
 sky130_fd_sc_hs__fill_2 FILLER_151_229 ();
 sky130_fd_sc_hs__fill_1 FILLER_151_231 ();
 sky130_fd_sc_hs__fill_2 FILLER_151_233 ();
 sky130_fd_sc_hs__fill_1 FILLER_151_235 ();
 sky130_fd_sc_hs__fill_4 FILLER_151_244 ();
 sky130_fd_sc_hs__fill_2 FILLER_151_248 ();
 sky130_fd_sc_hs__fill_4 FILLER_151_284 ();
 sky130_fd_sc_hs__fill_2 FILLER_151_288 ();
 sky130_fd_sc_hs__fill_8 FILLER_151_304 ();
 sky130_fd_sc_hs__fill_4 FILLER_151_312 ();
 sky130_fd_sc_hs__fill_1 FILLER_151_316 ();
 sky130_fd_sc_hs__fill_4 FILLER_151_325 ();
 sky130_fd_sc_hs__fill_1 FILLER_151_329 ();
 sky130_fd_sc_hs__fill_8 FILLER_151_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_151_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_151_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_151_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_151_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_151_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_151_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_151_405 ();
 sky130_fd_sc_hs__fill_4 FILLER_151_407 ();
 sky130_fd_sc_hs__fill_2 FILLER_151_411 ();
 sky130_fd_sc_hs__fill_1 FILLER_151_413 ();
 sky130_fd_sc_hs__fill_1 FILLER_151_417 ();
 sky130_fd_sc_hs__fill_8 FILLER_151_421 ();
 sky130_fd_sc_hs__fill_8 FILLER_151_429 ();
 sky130_fd_sc_hs__fill_8 FILLER_151_437 ();
 sky130_fd_sc_hs__fill_2 FILLER_151_451 ();
 sky130_fd_sc_hs__fill_1 FILLER_151_453 ();
 sky130_fd_sc_hs__fill_4 FILLER_151_457 ();
 sky130_fd_sc_hs__fill_2 FILLER_151_461 ();
 sky130_fd_sc_hs__fill_1 FILLER_151_463 ();
 sky130_fd_sc_hs__fill_2 FILLER_151_465 ();
 sky130_fd_sc_hs__fill_4 FILLER_151_518 ();
 sky130_fd_sc_hs__fill_1 FILLER_151_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_151_532 ();
 sky130_fd_sc_hs__fill_8 FILLER_152_0 ();
 sky130_fd_sc_hs__fill_2 FILLER_152_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_152_18 ();
 sky130_fd_sc_hs__fill_2 FILLER_152_26 ();
 sky130_fd_sc_hs__fill_1 FILLER_152_28 ();
 sky130_fd_sc_hs__fill_4 FILLER_152_30 ();
 sky130_fd_sc_hs__fill_1 FILLER_152_34 ();
 sky130_fd_sc_hs__fill_8 FILLER_152_75 ();
 sky130_fd_sc_hs__fill_4 FILLER_152_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_152_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_152_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_152_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_152_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_152_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_152_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_152_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_152_144 ();
 sky130_fd_sc_hs__fill_1 FILLER_152_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_152_150 ();
 sky130_fd_sc_hs__fill_8 FILLER_152_158 ();
 sky130_fd_sc_hs__fill_2 FILLER_152_166 ();
 sky130_fd_sc_hs__fill_2 FILLER_152_187 ();
 sky130_fd_sc_hs__fill_2 FILLER_152_196 ();
 sky130_fd_sc_hs__fill_1 FILLER_152_198 ();
 sky130_fd_sc_hs__fill_8 FILLER_152_219 ();
 sky130_fd_sc_hs__fill_4 FILLER_152_227 ();
 sky130_fd_sc_hs__fill_2 FILLER_152_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_152_247 ();
 sky130_fd_sc_hs__fill_4 FILLER_152_255 ();
 sky130_fd_sc_hs__fill_2 FILLER_152_259 ();
 sky130_fd_sc_hs__fill_8 FILLER_152_267 ();
 sky130_fd_sc_hs__fill_8 FILLER_152_275 ();
 sky130_fd_sc_hs__fill_2 FILLER_152_283 ();
 sky130_fd_sc_hs__fill_1 FILLER_152_285 ();
 sky130_fd_sc_hs__fill_8 FILLER_152_300 ();
 sky130_fd_sc_hs__fill_2 FILLER_152_308 ();
 sky130_fd_sc_hs__fill_4 FILLER_152_313 ();
 sky130_fd_sc_hs__fill_2 FILLER_152_317 ();
 sky130_fd_sc_hs__fill_8 FILLER_152_320 ();
 sky130_fd_sc_hs__fill_1 FILLER_152_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_152_350 ();
 sky130_fd_sc_hs__fill_8 FILLER_152_358 ();
 sky130_fd_sc_hs__fill_8 FILLER_152_366 ();
 sky130_fd_sc_hs__fill_2 FILLER_152_374 ();
 sky130_fd_sc_hs__fill_1 FILLER_152_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_152_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_152_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_152_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_152_402 ();
 sky130_fd_sc_hs__fill_1 FILLER_152_410 ();
 sky130_fd_sc_hs__fill_4 FILLER_152_430 ();
 sky130_fd_sc_hs__fill_1 FILLER_152_434 ();
 sky130_fd_sc_hs__fill_1 FILLER_152_436 ();
 sky130_fd_sc_hs__fill_1 FILLER_152_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_152_494 ();
 sky130_fd_sc_hs__fill_4 FILLER_152_502 ();
 sky130_fd_sc_hs__fill_2 FILLER_152_506 ();
 sky130_fd_sc_hs__fill_8 FILLER_152_512 ();
 sky130_fd_sc_hs__fill_4 FILLER_152_520 ();
 sky130_fd_sc_hs__fill_1 FILLER_152_524 ();
 sky130_fd_sc_hs__fill_4 FILLER_152_533 ();
 sky130_fd_sc_hs__fill_2 FILLER_152_537 ();
 sky130_fd_sc_hs__fill_1 FILLER_152_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_153_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_153_8 ();
 sky130_fd_sc_hs__fill_4 FILLER_153_16 ();
 sky130_fd_sc_hs__fill_1 FILLER_153_20 ();
 sky130_fd_sc_hs__fill_8 FILLER_153_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_153_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_153_56 ();
 sky130_fd_sc_hs__fill_1 FILLER_153_59 ();
 sky130_fd_sc_hs__fill_2 FILLER_153_64 ();
 sky130_fd_sc_hs__fill_1 FILLER_153_66 ();
 sky130_fd_sc_hs__fill_4 FILLER_153_81 ();
 sky130_fd_sc_hs__fill_2 FILLER_153_85 ();
 sky130_fd_sc_hs__fill_1 FILLER_153_87 ();
 sky130_fd_sc_hs__fill_8 FILLER_153_117 ();
 sky130_fd_sc_hs__fill_2 FILLER_153_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_153_156 ();
 sky130_fd_sc_hs__fill_8 FILLER_153_164 ();
 sky130_fd_sc_hs__fill_2 FILLER_153_172 ();
 sky130_fd_sc_hs__fill_8 FILLER_153_175 ();
 sky130_fd_sc_hs__fill_4 FILLER_153_183 ();
 sky130_fd_sc_hs__fill_1 FILLER_153_187 ();
 sky130_fd_sc_hs__fill_2 FILLER_153_195 ();
 sky130_fd_sc_hs__fill_1 FILLER_153_204 ();
 sky130_fd_sc_hs__fill_2 FILLER_153_209 ();
 sky130_fd_sc_hs__fill_8 FILLER_153_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_153_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_153_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_153_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_153_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_153_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_153_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_153_289 ();
 sky130_fd_sc_hs__fill_2 FILLER_153_299 ();
 sky130_fd_sc_hs__fill_1 FILLER_153_301 ();
 sky130_fd_sc_hs__fill_8 FILLER_153_319 ();
 sky130_fd_sc_hs__fill_8 FILLER_153_353 ();
 sky130_fd_sc_hs__fill_8 FILLER_153_361 ();
 sky130_fd_sc_hs__fill_4 FILLER_153_369 ();
 sky130_fd_sc_hs__fill_8 FILLER_153_423 ();
 sky130_fd_sc_hs__fill_4 FILLER_153_431 ();
 sky130_fd_sc_hs__fill_2 FILLER_153_435 ();
 sky130_fd_sc_hs__fill_4 FILLER_153_443 ();
 sky130_fd_sc_hs__fill_2 FILLER_153_447 ();
 sky130_fd_sc_hs__fill_1 FILLER_153_452 ();
 sky130_fd_sc_hs__fill_4 FILLER_153_457 ();
 sky130_fd_sc_hs__fill_2 FILLER_153_461 ();
 sky130_fd_sc_hs__fill_1 FILLER_153_463 ();
 sky130_fd_sc_hs__fill_2 FILLER_153_465 ();
 sky130_fd_sc_hs__fill_1 FILLER_153_467 ();
 sky130_fd_sc_hs__fill_4 FILLER_153_508 ();
 sky130_fd_sc_hs__fill_2 FILLER_153_512 ();
 sky130_fd_sc_hs__fill_8 FILLER_153_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_153_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_153_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_154_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_154_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_154_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_154_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_154_28 ();
 sky130_fd_sc_hs__fill_4 FILLER_154_30 ();
 sky130_fd_sc_hs__fill_1 FILLER_154_34 ();
 sky130_fd_sc_hs__fill_4 FILLER_154_69 ();
 sky130_fd_sc_hs__fill_2 FILLER_154_73 ();
 sky130_fd_sc_hs__fill_1 FILLER_154_75 ();
 sky130_fd_sc_hs__fill_4 FILLER_154_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_154_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_154_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_154_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_154_112 ();
 sky130_fd_sc_hs__fill_4 FILLER_154_120 ();
 sky130_fd_sc_hs__fill_1 FILLER_154_124 ();
 sky130_fd_sc_hs__fill_8 FILLER_154_132 ();
 sky130_fd_sc_hs__fill_4 FILLER_154_140 ();
 sky130_fd_sc_hs__fill_1 FILLER_154_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_154_146 ();
 sky130_fd_sc_hs__fill_4 FILLER_154_154 ();
 sky130_fd_sc_hs__fill_2 FILLER_154_158 ();
 sky130_fd_sc_hs__fill_1 FILLER_154_160 ();
 sky130_fd_sc_hs__fill_4 FILLER_154_168 ();
 sky130_fd_sc_hs__fill_2 FILLER_154_172 ();
 sky130_fd_sc_hs__fill_1 FILLER_154_174 ();
 sky130_fd_sc_hs__fill_4 FILLER_154_196 ();
 sky130_fd_sc_hs__fill_2 FILLER_154_200 ();
 sky130_fd_sc_hs__fill_1 FILLER_154_202 ();
 sky130_fd_sc_hs__fill_1 FILLER_154_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_154_208 ();
 sky130_fd_sc_hs__fill_8 FILLER_154_216 ();
 sky130_fd_sc_hs__fill_8 FILLER_154_224 ();
 sky130_fd_sc_hs__fill_8 FILLER_154_232 ();
 sky130_fd_sc_hs__fill_8 FILLER_154_240 ();
 sky130_fd_sc_hs__fill_4 FILLER_154_248 ();
 sky130_fd_sc_hs__fill_1 FILLER_154_252 ();
 sky130_fd_sc_hs__fill_8 FILLER_154_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_154_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_154_278 ();
 sky130_fd_sc_hs__fill_4 FILLER_154_286 ();
 sky130_fd_sc_hs__fill_2 FILLER_154_290 ();
 sky130_fd_sc_hs__fill_1 FILLER_154_292 ();
 sky130_fd_sc_hs__fill_8 FILLER_154_310 ();
 sky130_fd_sc_hs__fill_1 FILLER_154_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_154_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_154_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_154_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_154_344 ();
 sky130_fd_sc_hs__fill_4 FILLER_154_352 ();
 sky130_fd_sc_hs__fill_1 FILLER_154_356 ();
 sky130_fd_sc_hs__fill_2 FILLER_154_375 ();
 sky130_fd_sc_hs__fill_8 FILLER_154_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_154_386 ();
 sky130_fd_sc_hs__fill_4 FILLER_154_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_154_403 ();
 sky130_fd_sc_hs__fill_8 FILLER_154_411 ();
 sky130_fd_sc_hs__fill_2 FILLER_154_419 ();
 sky130_fd_sc_hs__fill_1 FILLER_154_421 ();
 sky130_fd_sc_hs__fill_8 FILLER_154_427 ();
 sky130_fd_sc_hs__fill_8 FILLER_154_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_154_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_154_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_154_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_154_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_154_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_154_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_154_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_154_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_154_502 ();
 sky130_fd_sc_hs__fill_2 FILLER_154_510 ();
 sky130_fd_sc_hs__fill_2 FILLER_154_515 ();
 sky130_fd_sc_hs__fill_8 FILLER_155_0 ();
 sky130_fd_sc_hs__fill_4 FILLER_155_8 ();
 sky130_fd_sc_hs__fill_2 FILLER_155_12 ();
 sky130_fd_sc_hs__fill_1 FILLER_155_14 ();
 sky130_fd_sc_hs__fill_8 FILLER_155_23 ();
 sky130_fd_sc_hs__fill_8 FILLER_155_31 ();
 sky130_fd_sc_hs__fill_8 FILLER_155_39 ();
 sky130_fd_sc_hs__fill_8 FILLER_155_47 ();
 sky130_fd_sc_hs__fill_2 FILLER_155_55 ();
 sky130_fd_sc_hs__fill_1 FILLER_155_57 ();
 sky130_fd_sc_hs__fill_8 FILLER_155_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_155_67 ();
 sky130_fd_sc_hs__fill_2 FILLER_155_75 ();
 sky130_fd_sc_hs__fill_1 FILLER_155_77 ();
 sky130_fd_sc_hs__fill_8 FILLER_155_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_155_94 ();
 sky130_fd_sc_hs__fill_4 FILLER_155_102 ();
 sky130_fd_sc_hs__fill_2 FILLER_155_106 ();
 sky130_fd_sc_hs__fill_2 FILLER_155_114 ();
 sky130_fd_sc_hs__fill_8 FILLER_155_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_155_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_155_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_155_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_155_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_155_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_155_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_155_173 ();
 sky130_fd_sc_hs__fill_1 FILLER_155_175 ();
 sky130_fd_sc_hs__fill_2 FILLER_155_180 ();
 sky130_fd_sc_hs__fill_8 FILLER_155_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_155_194 ();
 sky130_fd_sc_hs__fill_8 FILLER_155_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_155_210 ();
 sky130_fd_sc_hs__fill_8 FILLER_155_218 ();
 sky130_fd_sc_hs__fill_4 FILLER_155_226 ();
 sky130_fd_sc_hs__fill_2 FILLER_155_230 ();
 sky130_fd_sc_hs__fill_4 FILLER_155_233 ();
 sky130_fd_sc_hs__fill_1 FILLER_155_237 ();
 sky130_fd_sc_hs__fill_2 FILLER_155_245 ();
 sky130_fd_sc_hs__fill_1 FILLER_155_247 ();
 sky130_fd_sc_hs__fill_1 FILLER_155_280 ();
 sky130_fd_sc_hs__fill_4 FILLER_155_284 ();
 sky130_fd_sc_hs__fill_2 FILLER_155_288 ();
 sky130_fd_sc_hs__fill_8 FILLER_155_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_155_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_155_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_155_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_155_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_155_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_155_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_155_347 ();
 sky130_fd_sc_hs__fill_2 FILLER_155_349 ();
 sky130_fd_sc_hs__fill_1 FILLER_155_351 ();
 sky130_fd_sc_hs__fill_2 FILLER_155_373 ();
 sky130_fd_sc_hs__fill_1 FILLER_155_375 ();
 sky130_fd_sc_hs__fill_8 FILLER_155_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_155_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_155_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_155_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_155_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_155_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_155_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_155_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_155_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_155_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_155_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_155_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_155_481 ();
 sky130_fd_sc_hs__fill_2 FILLER_155_489 ();
 sky130_fd_sc_hs__fill_1 FILLER_155_491 ();
 sky130_fd_sc_hs__fill_8 FILLER_155_523 ();
 sky130_fd_sc_hs__fill_1 FILLER_155_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_156_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_156_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_156_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_156_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_156_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_156_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_156_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_156_54 ();
 sky130_fd_sc_hs__fill_4 FILLER_156_62 ();
 sky130_fd_sc_hs__fill_4 FILLER_156_81 ();
 sky130_fd_sc_hs__fill_2 FILLER_156_85 ();
 sky130_fd_sc_hs__fill_8 FILLER_156_88 ();
 sky130_fd_sc_hs__fill_1 FILLER_156_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_156_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_156_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_156_120 ();
 sky130_fd_sc_hs__fill_1 FILLER_156_128 ();
 sky130_fd_sc_hs__fill_2 FILLER_156_143 ();
 sky130_fd_sc_hs__fill_4 FILLER_156_146 ();
 sky130_fd_sc_hs__fill_2 FILLER_156_150 ();
 sky130_fd_sc_hs__fill_1 FILLER_156_152 ();
 sky130_fd_sc_hs__fill_2 FILLER_156_160 ();
 sky130_fd_sc_hs__fill_8 FILLER_156_165 ();
 sky130_fd_sc_hs__fill_8 FILLER_156_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_156_181 ();
 sky130_fd_sc_hs__fill_2 FILLER_156_189 ();
 sky130_fd_sc_hs__fill_8 FILLER_156_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_156_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_156_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_156_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_156_236 ();
 sky130_fd_sc_hs__fill_2 FILLER_156_244 ();
 sky130_fd_sc_hs__fill_1 FILLER_156_246 ();
 sky130_fd_sc_hs__fill_8 FILLER_156_262 ();
 sky130_fd_sc_hs__fill_2 FILLER_156_270 ();
 sky130_fd_sc_hs__fill_4 FILLER_156_289 ();
 sky130_fd_sc_hs__fill_1 FILLER_156_293 ();
 sky130_fd_sc_hs__fill_8 FILLER_156_303 ();
 sky130_fd_sc_hs__fill_8 FILLER_156_311 ();
 sky130_fd_sc_hs__fill_8 FILLER_156_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_156_328 ();
 sky130_fd_sc_hs__fill_4 FILLER_156_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_156_343 ();
 sky130_fd_sc_hs__fill_2 FILLER_156_351 ();
 sky130_fd_sc_hs__fill_1 FILLER_156_353 ();
 sky130_fd_sc_hs__fill_4 FILLER_156_371 ();
 sky130_fd_sc_hs__fill_2 FILLER_156_375 ();
 sky130_fd_sc_hs__fill_8 FILLER_156_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_156_386 ();
 sky130_fd_sc_hs__fill_4 FILLER_156_394 ();
 sky130_fd_sc_hs__fill_1 FILLER_156_398 ();
 sky130_fd_sc_hs__fill_8 FILLER_156_420 ();
 sky130_fd_sc_hs__fill_4 FILLER_156_428 ();
 sky130_fd_sc_hs__fill_2 FILLER_156_432 ();
 sky130_fd_sc_hs__fill_1 FILLER_156_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_156_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_156_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_156_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_156_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_156_468 ();
 sky130_fd_sc_hs__fill_2 FILLER_156_476 ();
 sky130_fd_sc_hs__fill_1 FILLER_156_478 ();
 sky130_fd_sc_hs__fill_8 FILLER_156_494 ();
 sky130_fd_sc_hs__fill_4 FILLER_156_502 ();
 sky130_fd_sc_hs__fill_2 FILLER_156_506 ();
 sky130_fd_sc_hs__fill_1 FILLER_156_508 ();
 sky130_fd_sc_hs__fill_1 FILLER_156_516 ();
 sky130_fd_sc_hs__fill_8 FILLER_157_0 ();
 sky130_fd_sc_hs__fill_4 FILLER_157_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_157_20 ();
 sky130_fd_sc_hs__fill_8 FILLER_157_28 ();
 sky130_fd_sc_hs__fill_2 FILLER_157_36 ();
 sky130_fd_sc_hs__fill_1 FILLER_157_38 ();
 sky130_fd_sc_hs__fill_1 FILLER_157_57 ();
 sky130_fd_sc_hs__fill_8 FILLER_157_59 ();
 sky130_fd_sc_hs__fill_1 FILLER_157_67 ();
 sky130_fd_sc_hs__fill_2 FILLER_157_76 ();
 sky130_fd_sc_hs__fill_8 FILLER_157_93 ();
 sky130_fd_sc_hs__fill_1 FILLER_157_101 ();
 sky130_fd_sc_hs__fill_1 FILLER_157_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_157_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_157_125 ();
 sky130_fd_sc_hs__fill_1 FILLER_157_139 ();
 sky130_fd_sc_hs__fill_4 FILLER_157_146 ();
 sky130_fd_sc_hs__fill_2 FILLER_157_171 ();
 sky130_fd_sc_hs__fill_1 FILLER_157_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_157_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_157_183 ();
 sky130_fd_sc_hs__fill_2 FILLER_157_191 ();
 sky130_fd_sc_hs__fill_1 FILLER_157_193 ();
 sky130_fd_sc_hs__fill_1 FILLER_157_201 ();
 sky130_fd_sc_hs__fill_8 FILLER_157_217 ();
 sky130_fd_sc_hs__fill_4 FILLER_157_225 ();
 sky130_fd_sc_hs__fill_2 FILLER_157_229 ();
 sky130_fd_sc_hs__fill_1 FILLER_157_231 ();
 sky130_fd_sc_hs__fill_4 FILLER_157_233 ();
 sky130_fd_sc_hs__fill_1 FILLER_157_237 ();
 sky130_fd_sc_hs__fill_1 FILLER_157_254 ();
 sky130_fd_sc_hs__fill_1 FILLER_157_258 ();
 sky130_fd_sc_hs__fill_2 FILLER_157_263 ();
 sky130_fd_sc_hs__fill_2 FILLER_157_291 ();
 sky130_fd_sc_hs__fill_1 FILLER_157_293 ();
 sky130_fd_sc_hs__fill_8 FILLER_157_301 ();
 sky130_fd_sc_hs__fill_1 FILLER_157_309 ();
 sky130_fd_sc_hs__fill_8 FILLER_157_313 ();
 sky130_fd_sc_hs__fill_8 FILLER_157_321 ();
 sky130_fd_sc_hs__fill_2 FILLER_157_329 ();
 sky130_fd_sc_hs__fill_1 FILLER_157_331 ();
 sky130_fd_sc_hs__fill_2 FILLER_157_345 ();
 sky130_fd_sc_hs__fill_1 FILLER_157_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_157_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_157_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_157_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_157_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_157_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_157_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_157_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_157_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_157_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_157_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_157_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_157_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_157_439 ();
 sky130_fd_sc_hs__fill_4 FILLER_157_447 ();
 sky130_fd_sc_hs__fill_2 FILLER_157_461 ();
 sky130_fd_sc_hs__fill_1 FILLER_157_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_157_493 ();
 sky130_fd_sc_hs__fill_2 FILLER_157_501 ();
 sky130_fd_sc_hs__fill_1 FILLER_157_503 ();
 sky130_fd_sc_hs__fill_1 FILLER_157_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_158_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_158_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_158_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_158_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_158_28 ();
 sky130_fd_sc_hs__fill_4 FILLER_158_30 ();
 sky130_fd_sc_hs__fill_1 FILLER_158_34 ();
 sky130_fd_sc_hs__fill_2 FILLER_158_42 ();
 sky130_fd_sc_hs__fill_1 FILLER_158_44 ();
 sky130_fd_sc_hs__fill_2 FILLER_158_64 ();
 sky130_fd_sc_hs__fill_1 FILLER_158_66 ();
 sky130_fd_sc_hs__fill_4 FILLER_158_82 ();
 sky130_fd_sc_hs__fill_1 FILLER_158_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_158_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_158_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_158_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_158_112 ();
 sky130_fd_sc_hs__fill_2 FILLER_158_128 ();
 sky130_fd_sc_hs__fill_4 FILLER_158_146 ();
 sky130_fd_sc_hs__fill_4 FILLER_158_166 ();
 sky130_fd_sc_hs__fill_2 FILLER_158_170 ();
 sky130_fd_sc_hs__fill_1 FILLER_158_172 ();
 sky130_fd_sc_hs__fill_8 FILLER_158_177 ();
 sky130_fd_sc_hs__fill_2 FILLER_158_185 ();
 sky130_fd_sc_hs__fill_1 FILLER_158_187 ();
 sky130_fd_sc_hs__fill_8 FILLER_158_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_158_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_158_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_158_228 ();
 sky130_fd_sc_hs__fill_2 FILLER_158_236 ();
 sky130_fd_sc_hs__fill_1 FILLER_158_238 ();
 sky130_fd_sc_hs__fill_4 FILLER_158_254 ();
 sky130_fd_sc_hs__fill_2 FILLER_158_258 ();
 sky130_fd_sc_hs__fill_1 FILLER_158_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_158_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_158_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_158_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_158_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_158_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_158_320 ();
 sky130_fd_sc_hs__fill_4 FILLER_158_328 ();
 sky130_fd_sc_hs__fill_1 FILLER_158_332 ();
 sky130_fd_sc_hs__fill_4 FILLER_158_372 ();
 sky130_fd_sc_hs__fill_1 FILLER_158_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_158_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_158_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_158_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_158_402 ();
 sky130_fd_sc_hs__fill_2 FILLER_158_410 ();
 sky130_fd_sc_hs__fill_1 FILLER_158_412 ();
 sky130_fd_sc_hs__fill_8 FILLER_158_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_158_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_158_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_158_470 ();
 sky130_fd_sc_hs__fill_8 FILLER_158_478 ();
 sky130_fd_sc_hs__fill_4 FILLER_158_486 ();
 sky130_fd_sc_hs__fill_2 FILLER_158_490 ();
 sky130_fd_sc_hs__fill_1 FILLER_158_492 ();
 sky130_fd_sc_hs__fill_4 FILLER_158_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_158_505 ();
 sky130_fd_sc_hs__fill_1 FILLER_158_513 ();
 sky130_fd_sc_hs__fill_8 FILLER_158_522 ();
 sky130_fd_sc_hs__fill_8 FILLER_158_530 ();
 sky130_fd_sc_hs__fill_2 FILLER_158_538 ();
 sky130_fd_sc_hs__fill_4 FILLER_159_0 ();
 sky130_fd_sc_hs__fill_2 FILLER_159_4 ();
 sky130_fd_sc_hs__fill_1 FILLER_159_6 ();
 sky130_fd_sc_hs__fill_4 FILLER_159_33 ();
 sky130_fd_sc_hs__fill_2 FILLER_159_59 ();
 sky130_fd_sc_hs__fill_1 FILLER_159_61 ();
 sky130_fd_sc_hs__fill_8 FILLER_159_66 ();
 sky130_fd_sc_hs__fill_8 FILLER_159_74 ();
 sky130_fd_sc_hs__fill_8 FILLER_159_82 ();
 sky130_fd_sc_hs__fill_8 FILLER_159_90 ();
 sky130_fd_sc_hs__fill_8 FILLER_159_98 ();
 sky130_fd_sc_hs__fill_8 FILLER_159_106 ();
 sky130_fd_sc_hs__fill_2 FILLER_159_114 ();
 sky130_fd_sc_hs__fill_4 FILLER_159_117 ();
 sky130_fd_sc_hs__fill_2 FILLER_159_121 ();
 sky130_fd_sc_hs__fill_1 FILLER_159_123 ();
 sky130_fd_sc_hs__fill_4 FILLER_159_168 ();
 sky130_fd_sc_hs__fill_2 FILLER_159_172 ();
 sky130_fd_sc_hs__fill_8 FILLER_159_175 ();
 sky130_fd_sc_hs__fill_4 FILLER_159_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_159_195 ();
 sky130_fd_sc_hs__fill_8 FILLER_159_203 ();
 sky130_fd_sc_hs__fill_8 FILLER_159_211 ();
 sky130_fd_sc_hs__fill_8 FILLER_159_219 ();
 sky130_fd_sc_hs__fill_4 FILLER_159_227 ();
 sky130_fd_sc_hs__fill_1 FILLER_159_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_159_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_159_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_159_249 ();
 sky130_fd_sc_hs__fill_4 FILLER_159_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_159_269 ();
 sky130_fd_sc_hs__fill_8 FILLER_159_277 ();
 sky130_fd_sc_hs__fill_4 FILLER_159_285 ();
 sky130_fd_sc_hs__fill_1 FILLER_159_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_159_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_159_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_159_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_159_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_159_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_159_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_159_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_159_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_159_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_159_357 ();
 sky130_fd_sc_hs__fill_2 FILLER_159_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_159_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_159_384 ();
 sky130_fd_sc_hs__fill_8 FILLER_159_392 ();
 sky130_fd_sc_hs__fill_4 FILLER_159_400 ();
 sky130_fd_sc_hs__fill_2 FILLER_159_404 ();
 sky130_fd_sc_hs__fill_2 FILLER_159_407 ();
 sky130_fd_sc_hs__fill_1 FILLER_159_409 ();
 sky130_fd_sc_hs__fill_8 FILLER_159_414 ();
 sky130_fd_sc_hs__fill_8 FILLER_159_422 ();
 sky130_fd_sc_hs__fill_8 FILLER_159_430 ();
 sky130_fd_sc_hs__fill_8 FILLER_159_438 ();
 sky130_fd_sc_hs__fill_8 FILLER_159_446 ();
 sky130_fd_sc_hs__fill_4 FILLER_159_454 ();
 sky130_fd_sc_hs__fill_8 FILLER_159_465 ();
 sky130_fd_sc_hs__fill_2 FILLER_159_473 ();
 sky130_fd_sc_hs__fill_1 FILLER_159_475 ();
 sky130_fd_sc_hs__fill_8 FILLER_159_494 ();
 sky130_fd_sc_hs__fill_1 FILLER_159_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_159_506 ();
 sky130_fd_sc_hs__fill_8 FILLER_159_514 ();
 sky130_fd_sc_hs__fill_8 FILLER_159_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_159_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_159_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_160_0 ();
 sky130_fd_sc_hs__fill_2 FILLER_160_8 ();
 sky130_fd_sc_hs__fill_1 FILLER_160_18 ();
 sky130_fd_sc_hs__fill_2 FILLER_160_30 ();
 sky130_fd_sc_hs__fill_1 FILLER_160_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_160_46 ();
 sky130_fd_sc_hs__fill_4 FILLER_160_54 ();
 sky130_fd_sc_hs__fill_2 FILLER_160_58 ();
 sky130_fd_sc_hs__fill_1 FILLER_160_60 ();
 sky130_fd_sc_hs__fill_8 FILLER_160_74 ();
 sky130_fd_sc_hs__fill_4 FILLER_160_82 ();
 sky130_fd_sc_hs__fill_1 FILLER_160_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_160_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_160_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_160_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_160_112 ();
 sky130_fd_sc_hs__fill_2 FILLER_160_120 ();
 sky130_fd_sc_hs__fill_1 FILLER_160_122 ();
 sky130_fd_sc_hs__fill_8 FILLER_160_131 ();
 sky130_fd_sc_hs__fill_4 FILLER_160_139 ();
 sky130_fd_sc_hs__fill_2 FILLER_160_143 ();
 sky130_fd_sc_hs__fill_4 FILLER_160_153 ();
 sky130_fd_sc_hs__fill_1 FILLER_160_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_160_165 ();
 sky130_fd_sc_hs__fill_8 FILLER_160_173 ();
 sky130_fd_sc_hs__fill_2 FILLER_160_181 ();
 sky130_fd_sc_hs__fill_1 FILLER_160_183 ();
 sky130_fd_sc_hs__fill_2 FILLER_160_192 ();
 sky130_fd_sc_hs__fill_1 FILLER_160_194 ();
 sky130_fd_sc_hs__fill_8 FILLER_160_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_160_212 ();
 sky130_fd_sc_hs__fill_4 FILLER_160_220 ();
 sky130_fd_sc_hs__fill_2 FILLER_160_238 ();
 sky130_fd_sc_hs__fill_8 FILLER_160_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_160_260 ();
 sky130_fd_sc_hs__fill_2 FILLER_160_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_160_267 ();
 sky130_fd_sc_hs__fill_8 FILLER_160_275 ();
 sky130_fd_sc_hs__fill_8 FILLER_160_283 ();
 sky130_fd_sc_hs__fill_8 FILLER_160_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_160_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_160_307 ();
 sky130_fd_sc_hs__fill_4 FILLER_160_315 ();
 sky130_fd_sc_hs__fill_2 FILLER_160_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_160_335 ();
 sky130_fd_sc_hs__fill_4 FILLER_160_343 ();
 sky130_fd_sc_hs__fill_2 FILLER_160_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_160_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_160_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_160_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_160_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_160_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_160_386 ();
 sky130_fd_sc_hs__fill_4 FILLER_160_394 ();
 sky130_fd_sc_hs__fill_2 FILLER_160_398 ();
 sky130_fd_sc_hs__fill_8 FILLER_160_417 ();
 sky130_fd_sc_hs__fill_8 FILLER_160_425 ();
 sky130_fd_sc_hs__fill_2 FILLER_160_433 ();
 sky130_fd_sc_hs__fill_8 FILLER_160_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_160_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_160_452 ();
 sky130_fd_sc_hs__fill_2 FILLER_160_460 ();
 sky130_fd_sc_hs__fill_1 FILLER_160_468 ();
 sky130_fd_sc_hs__fill_4 FILLER_160_486 ();
 sky130_fd_sc_hs__fill_2 FILLER_160_490 ();
 sky130_fd_sc_hs__fill_1 FILLER_160_492 ();
 sky130_fd_sc_hs__fill_4 FILLER_160_494 ();
 sky130_fd_sc_hs__fill_2 FILLER_160_509 ();
 sky130_fd_sc_hs__fill_1 FILLER_160_511 ();
 sky130_fd_sc_hs__fill_4 FILLER_161_0 ();
 sky130_fd_sc_hs__fill_2 FILLER_161_4 ();
 sky130_fd_sc_hs__fill_1 FILLER_161_6 ();
 sky130_fd_sc_hs__fill_8 FILLER_161_15 ();
 sky130_fd_sc_hs__fill_8 FILLER_161_26 ();
 sky130_fd_sc_hs__fill_2 FILLER_161_34 ();
 sky130_fd_sc_hs__fill_4 FILLER_161_51 ();
 sky130_fd_sc_hs__fill_2 FILLER_161_55 ();
 sky130_fd_sc_hs__fill_1 FILLER_161_57 ();
 sky130_fd_sc_hs__fill_8 FILLER_161_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_161_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_161_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_161_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_161_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_161_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_161_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_161_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_161_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_161_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_161_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_161_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_161_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_161_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_161_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_161_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_161_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_161_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_161_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_161_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_161_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_161_215 ();
 sky130_fd_sc_hs__fill_2 FILLER_161_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_161_250 ();
 sky130_fd_sc_hs__fill_8 FILLER_161_258 ();
 sky130_fd_sc_hs__fill_8 FILLER_161_270 ();
 sky130_fd_sc_hs__fill_2 FILLER_161_278 ();
 sky130_fd_sc_hs__fill_1 FILLER_161_280 ();
 sky130_fd_sc_hs__fill_4 FILLER_161_284 ();
 sky130_fd_sc_hs__fill_2 FILLER_161_288 ();
 sky130_fd_sc_hs__fill_8 FILLER_161_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_161_299 ();
 sky130_fd_sc_hs__fill_4 FILLER_161_307 ();
 sky130_fd_sc_hs__fill_4 FILLER_161_320 ();
 sky130_fd_sc_hs__fill_2 FILLER_161_324 ();
 sky130_fd_sc_hs__fill_1 FILLER_161_326 ();
 sky130_fd_sc_hs__fill_4 FILLER_161_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_161_354 ();
 sky130_fd_sc_hs__fill_8 FILLER_161_362 ();
 sky130_fd_sc_hs__fill_8 FILLER_161_370 ();
 sky130_fd_sc_hs__fill_8 FILLER_161_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_161_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_161_394 ();
 sky130_fd_sc_hs__fill_4 FILLER_161_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_161_414 ();
 sky130_fd_sc_hs__fill_8 FILLER_161_422 ();
 sky130_fd_sc_hs__fill_8 FILLER_161_430 ();
 sky130_fd_sc_hs__fill_4 FILLER_161_438 ();
 sky130_fd_sc_hs__fill_8 FILLER_161_448 ();
 sky130_fd_sc_hs__fill_8 FILLER_161_456 ();
 sky130_fd_sc_hs__fill_8 FILLER_161_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_161_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_161_481 ();
 sky130_fd_sc_hs__fill_1 FILLER_161_489 ();
 sky130_fd_sc_hs__fill_2 FILLER_161_519 ();
 sky130_fd_sc_hs__fill_1 FILLER_161_521 ();
 sky130_fd_sc_hs__fill_1 FILLER_161_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_161_532 ();
 sky130_fd_sc_hs__fill_8 FILLER_162_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_162_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_162_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_162_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_162_28 ();
 sky130_fd_sc_hs__fill_4 FILLER_162_53 ();
 sky130_fd_sc_hs__fill_8 FILLER_162_64 ();
 sky130_fd_sc_hs__fill_4 FILLER_162_72 ();
 sky130_fd_sc_hs__fill_4 FILLER_162_88 ();
 sky130_fd_sc_hs__fill_2 FILLER_162_92 ();
 sky130_fd_sc_hs__fill_8 FILLER_162_113 ();
 sky130_fd_sc_hs__fill_8 FILLER_162_121 ();
 sky130_fd_sc_hs__fill_8 FILLER_162_129 ();
 sky130_fd_sc_hs__fill_8 FILLER_162_137 ();
 sky130_fd_sc_hs__fill_8 FILLER_162_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_162_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_162_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_162_170 ();
 sky130_fd_sc_hs__fill_4 FILLER_162_178 ();
 sky130_fd_sc_hs__fill_2 FILLER_162_182 ();
 sky130_fd_sc_hs__fill_8 FILLER_162_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_162_212 ();
 sky130_fd_sc_hs__fill_2 FILLER_162_220 ();
 sky130_fd_sc_hs__fill_1 FILLER_162_222 ();
 sky130_fd_sc_hs__fill_8 FILLER_162_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_162_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_162_260 ();
 sky130_fd_sc_hs__fill_4 FILLER_162_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_162_281 ();
 sky130_fd_sc_hs__fill_8 FILLER_162_289 ();
 sky130_fd_sc_hs__fill_2 FILLER_162_297 ();
 sky130_fd_sc_hs__fill_1 FILLER_162_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_162_308 ();
 sky130_fd_sc_hs__fill_2 FILLER_162_316 ();
 sky130_fd_sc_hs__fill_1 FILLER_162_318 ();
 sky130_fd_sc_hs__fill_4 FILLER_162_320 ();
 sky130_fd_sc_hs__fill_1 FILLER_162_339 ();
 sky130_fd_sc_hs__fill_8 FILLER_162_345 ();
 sky130_fd_sc_hs__fill_8 FILLER_162_353 ();
 sky130_fd_sc_hs__fill_2 FILLER_162_361 ();
 sky130_fd_sc_hs__fill_1 FILLER_162_363 ();
 sky130_fd_sc_hs__fill_8 FILLER_162_369 ();
 sky130_fd_sc_hs__fill_8 FILLER_162_378 ();
 sky130_fd_sc_hs__fill_2 FILLER_162_386 ();
 sky130_fd_sc_hs__fill_1 FILLER_162_388 ();
 sky130_fd_sc_hs__fill_8 FILLER_162_398 ();
 sky130_fd_sc_hs__fill_2 FILLER_162_406 ();
 sky130_fd_sc_hs__fill_8 FILLER_162_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_162_423 ();
 sky130_fd_sc_hs__fill_4 FILLER_162_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_162_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_162_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_162_452 ();
 sky130_fd_sc_hs__fill_2 FILLER_162_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_162_474 ();
 sky130_fd_sc_hs__fill_8 FILLER_162_482 ();
 sky130_fd_sc_hs__fill_2 FILLER_162_490 ();
 sky130_fd_sc_hs__fill_1 FILLER_162_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_162_494 ();
 sky130_fd_sc_hs__fill_4 FILLER_162_502 ();
 sky130_fd_sc_hs__fill_2 FILLER_162_506 ();
 sky130_fd_sc_hs__fill_1 FILLER_162_508 ();
 sky130_fd_sc_hs__fill_4 FILLER_162_535 ();
 sky130_fd_sc_hs__fill_1 FILLER_162_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_163_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_163_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_163_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_163_24 ();
 sky130_fd_sc_hs__fill_2 FILLER_163_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_163_41 ();
 sky130_fd_sc_hs__fill_8 FILLER_163_49 ();
 sky130_fd_sc_hs__fill_1 FILLER_163_57 ();
 sky130_fd_sc_hs__fill_8 FILLER_163_59 ();
 sky130_fd_sc_hs__fill_1 FILLER_163_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_163_106 ();
 sky130_fd_sc_hs__fill_2 FILLER_163_114 ();
 sky130_fd_sc_hs__fill_8 FILLER_163_117 ();
 sky130_fd_sc_hs__fill_1 FILLER_163_154 ();
 sky130_fd_sc_hs__fill_4 FILLER_163_175 ();
 sky130_fd_sc_hs__fill_2 FILLER_163_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_163_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_163_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_163_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_163_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_163_233 ();
 sky130_fd_sc_hs__fill_1 FILLER_163_241 ();
 sky130_fd_sc_hs__fill_1 FILLER_163_262 ();
 sky130_fd_sc_hs__fill_1 FILLER_163_271 ();
 sky130_fd_sc_hs__fill_1 FILLER_163_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_163_291 ();
 sky130_fd_sc_hs__fill_1 FILLER_163_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_163_303 ();
 sky130_fd_sc_hs__fill_8 FILLER_163_311 ();
 sky130_fd_sc_hs__fill_8 FILLER_163_319 ();
 sky130_fd_sc_hs__fill_4 FILLER_163_349 ();
 sky130_fd_sc_hs__fill_4 FILLER_163_360 ();
 sky130_fd_sc_hs__fill_4 FILLER_163_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_163_372 ();
 sky130_fd_sc_hs__fill_4 FILLER_163_380 ();
 sky130_fd_sc_hs__fill_1 FILLER_163_384 ();
 sky130_fd_sc_hs__fill_8 FILLER_163_391 ();
 sky130_fd_sc_hs__fill_4 FILLER_163_399 ();
 sky130_fd_sc_hs__fill_2 FILLER_163_403 ();
 sky130_fd_sc_hs__fill_1 FILLER_163_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_163_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_163_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_163_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_163_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_163_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_163_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_163_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_163_463 ();
 sky130_fd_sc_hs__fill_4 FILLER_163_465 ();
 sky130_fd_sc_hs__fill_2 FILLER_163_469 ();
 sky130_fd_sc_hs__fill_1 FILLER_163_471 ();
 sky130_fd_sc_hs__fill_8 FILLER_163_485 ();
 sky130_fd_sc_hs__fill_4 FILLER_163_493 ();
 sky130_fd_sc_hs__fill_1 FILLER_163_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_163_506 ();
 sky130_fd_sc_hs__fill_8 FILLER_163_514 ();
 sky130_fd_sc_hs__fill_2 FILLER_163_523 ();
 sky130_fd_sc_hs__fill_4 FILLER_163_533 ();
 sky130_fd_sc_hs__fill_2 FILLER_163_537 ();
 sky130_fd_sc_hs__fill_1 FILLER_163_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_164_8 ();
 sky130_fd_sc_hs__fill_4 FILLER_164_16 ();
 sky130_fd_sc_hs__fill_1 FILLER_164_20 ();
 sky130_fd_sc_hs__fill_8 FILLER_164_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_164_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_164_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_164_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_164_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_164_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_164_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_164_86 ();
 sky130_fd_sc_hs__fill_4 FILLER_164_88 ();
 sky130_fd_sc_hs__fill_2 FILLER_164_92 ();
 sky130_fd_sc_hs__fill_8 FILLER_164_105 ();
 sky130_fd_sc_hs__fill_8 FILLER_164_113 ();
 sky130_fd_sc_hs__fill_1 FILLER_164_121 ();
 sky130_fd_sc_hs__fill_4 FILLER_164_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_164_146 ();
 sky130_fd_sc_hs__fill_2 FILLER_164_154 ();
 sky130_fd_sc_hs__fill_1 FILLER_164_156 ();
 sky130_fd_sc_hs__fill_8 FILLER_164_164 ();
 sky130_fd_sc_hs__fill_4 FILLER_164_172 ();
 sky130_fd_sc_hs__fill_2 FILLER_164_176 ();
 sky130_fd_sc_hs__fill_8 FILLER_164_185 ();
 sky130_fd_sc_hs__fill_8 FILLER_164_193 ();
 sky130_fd_sc_hs__fill_2 FILLER_164_201 ();
 sky130_fd_sc_hs__fill_8 FILLER_164_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_164_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_164_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_164_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_164_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_164_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_164_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_164_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_164_262 ();
 sky130_fd_sc_hs__fill_4 FILLER_164_273 ();
 sky130_fd_sc_hs__fill_2 FILLER_164_277 ();
 sky130_fd_sc_hs__fill_4 FILLER_164_287 ();
 sky130_fd_sc_hs__fill_1 FILLER_164_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_164_309 ();
 sky130_fd_sc_hs__fill_2 FILLER_164_317 ();
 sky130_fd_sc_hs__fill_8 FILLER_164_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_164_328 ();
 sky130_fd_sc_hs__fill_2 FILLER_164_336 ();
 sky130_fd_sc_hs__fill_2 FILLER_164_355 ();
 sky130_fd_sc_hs__fill_1 FILLER_164_357 ();
 sky130_fd_sc_hs__fill_4 FILLER_164_370 ();
 sky130_fd_sc_hs__fill_2 FILLER_164_374 ();
 sky130_fd_sc_hs__fill_1 FILLER_164_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_164_378 ();
 sky130_fd_sc_hs__fill_4 FILLER_164_386 ();
 sky130_fd_sc_hs__fill_2 FILLER_164_390 ();
 sky130_fd_sc_hs__fill_1 FILLER_164_392 ();
 sky130_fd_sc_hs__fill_8 FILLER_164_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_164_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_164_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_164_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_164_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_164_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_164_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_164_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_164_460 ();
 sky130_fd_sc_hs__fill_4 FILLER_164_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_164_498 ();
 sky130_fd_sc_hs__fill_8 FILLER_164_506 ();
 sky130_fd_sc_hs__fill_8 FILLER_164_514 ();
 sky130_fd_sc_hs__fill_8 FILLER_164_522 ();
 sky130_fd_sc_hs__fill_8 FILLER_164_530 ();
 sky130_fd_sc_hs__fill_2 FILLER_164_538 ();
 sky130_fd_sc_hs__fill_8 FILLER_165_0 ();
 sky130_fd_sc_hs__fill_2 FILLER_165_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_165_18 ();
 sky130_fd_sc_hs__fill_1 FILLER_165_26 ();
 sky130_fd_sc_hs__fill_8 FILLER_165_44 ();
 sky130_fd_sc_hs__fill_4 FILLER_165_52 ();
 sky130_fd_sc_hs__fill_2 FILLER_165_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_165_59 ();
 sky130_fd_sc_hs__fill_1 FILLER_165_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_165_79 ();
 sky130_fd_sc_hs__fill_4 FILLER_165_87 ();
 sky130_fd_sc_hs__fill_2 FILLER_165_91 ();
 sky130_fd_sc_hs__fill_4 FILLER_165_112 ();
 sky130_fd_sc_hs__fill_1 FILLER_165_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_165_129 ();
 sky130_fd_sc_hs__fill_4 FILLER_165_137 ();
 sky130_fd_sc_hs__fill_8 FILLER_165_148 ();
 sky130_fd_sc_hs__fill_8 FILLER_165_156 ();
 sky130_fd_sc_hs__fill_8 FILLER_165_164 ();
 sky130_fd_sc_hs__fill_2 FILLER_165_172 ();
 sky130_fd_sc_hs__fill_8 FILLER_165_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_165_190 ();
 sky130_fd_sc_hs__fill_8 FILLER_165_198 ();
 sky130_fd_sc_hs__fill_8 FILLER_165_219 ();
 sky130_fd_sc_hs__fill_4 FILLER_165_227 ();
 sky130_fd_sc_hs__fill_1 FILLER_165_231 ();
 sky130_fd_sc_hs__fill_4 FILLER_165_233 ();
 sky130_fd_sc_hs__fill_1 FILLER_165_237 ();
 sky130_fd_sc_hs__fill_8 FILLER_165_243 ();
 sky130_fd_sc_hs__fill_8 FILLER_165_251 ();
 sky130_fd_sc_hs__fill_8 FILLER_165_259 ();
 sky130_fd_sc_hs__fill_8 FILLER_165_275 ();
 sky130_fd_sc_hs__fill_4 FILLER_165_283 ();
 sky130_fd_sc_hs__fill_8 FILLER_165_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_165_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_165_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_165_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_165_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_165_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_165_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_165_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_165_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_165_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_165_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_165_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_165_381 ();
 sky130_fd_sc_hs__fill_4 FILLER_165_389 ();
 sky130_fd_sc_hs__fill_2 FILLER_165_393 ();
 sky130_fd_sc_hs__fill_8 FILLER_165_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_165_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_165_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_165_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_165_439 ();
 sky130_fd_sc_hs__fill_4 FILLER_165_447 ();
 sky130_fd_sc_hs__fill_2 FILLER_165_451 ();
 sky130_fd_sc_hs__fill_1 FILLER_165_453 ();
 sky130_fd_sc_hs__fill_2 FILLER_165_461 ();
 sky130_fd_sc_hs__fill_1 FILLER_165_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_165_465 ();
 sky130_fd_sc_hs__fill_4 FILLER_165_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_165_503 ();
 sky130_fd_sc_hs__fill_8 FILLER_165_511 ();
 sky130_fd_sc_hs__fill_2 FILLER_165_519 ();
 sky130_fd_sc_hs__fill_1 FILLER_165_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_165_523 ();
 sky130_fd_sc_hs__fill_1 FILLER_165_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_166_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_166_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_166_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_166_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_166_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_166_30 ();
 sky130_fd_sc_hs__fill_4 FILLER_166_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_166_64 ();
 sky130_fd_sc_hs__fill_8 FILLER_166_72 ();
 sky130_fd_sc_hs__fill_4 FILLER_166_80 ();
 sky130_fd_sc_hs__fill_2 FILLER_166_84 ();
 sky130_fd_sc_hs__fill_1 FILLER_166_86 ();
 sky130_fd_sc_hs__fill_2 FILLER_166_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_166_112 ();
 sky130_fd_sc_hs__fill_4 FILLER_166_120 ();
 sky130_fd_sc_hs__fill_2 FILLER_166_124 ();
 sky130_fd_sc_hs__fill_1 FILLER_166_126 ();
 sky130_fd_sc_hs__fill_4 FILLER_166_139 ();
 sky130_fd_sc_hs__fill_2 FILLER_166_143 ();
 sky130_fd_sc_hs__fill_4 FILLER_166_146 ();
 sky130_fd_sc_hs__fill_2 FILLER_166_150 ();
 sky130_fd_sc_hs__fill_1 FILLER_166_152 ();
 sky130_fd_sc_hs__fill_2 FILLER_166_172 ();
 sky130_fd_sc_hs__fill_2 FILLER_166_181 ();
 sky130_fd_sc_hs__fill_1 FILLER_166_183 ();
 sky130_fd_sc_hs__fill_2 FILLER_166_204 ();
 sky130_fd_sc_hs__fill_1 FILLER_166_206 ();
 sky130_fd_sc_hs__fill_8 FILLER_166_225 ();
 sky130_fd_sc_hs__fill_8 FILLER_166_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_166_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_166_249 ();
 sky130_fd_sc_hs__fill_4 FILLER_166_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_166_280 ();
 sky130_fd_sc_hs__fill_8 FILLER_166_288 ();
 sky130_fd_sc_hs__fill_8 FILLER_166_296 ();
 sky130_fd_sc_hs__fill_8 FILLER_166_304 ();
 sky130_fd_sc_hs__fill_4 FILLER_166_312 ();
 sky130_fd_sc_hs__fill_2 FILLER_166_316 ();
 sky130_fd_sc_hs__fill_1 FILLER_166_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_166_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_166_334 ();
 sky130_fd_sc_hs__fill_8 FILLER_166_342 ();
 sky130_fd_sc_hs__fill_8 FILLER_166_350 ();
 sky130_fd_sc_hs__fill_8 FILLER_166_358 ();
 sky130_fd_sc_hs__fill_8 FILLER_166_366 ();
 sky130_fd_sc_hs__fill_2 FILLER_166_374 ();
 sky130_fd_sc_hs__fill_1 FILLER_166_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_166_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_166_386 ();
 sky130_fd_sc_hs__fill_4 FILLER_166_394 ();
 sky130_fd_sc_hs__fill_2 FILLER_166_398 ();
 sky130_fd_sc_hs__fill_8 FILLER_166_417 ();
 sky130_fd_sc_hs__fill_8 FILLER_166_425 ();
 sky130_fd_sc_hs__fill_2 FILLER_166_433 ();
 sky130_fd_sc_hs__fill_8 FILLER_166_436 ();
 sky130_fd_sc_hs__fill_2 FILLER_166_444 ();
 sky130_fd_sc_hs__fill_1 FILLER_166_446 ();
 sky130_fd_sc_hs__fill_8 FILLER_166_470 ();
 sky130_fd_sc_hs__fill_8 FILLER_166_478 ();
 sky130_fd_sc_hs__fill_4 FILLER_166_486 ();
 sky130_fd_sc_hs__fill_1 FILLER_166_494 ();
 sky130_fd_sc_hs__fill_4 FILLER_166_499 ();
 sky130_fd_sc_hs__fill_2 FILLER_166_503 ();
 sky130_fd_sc_hs__fill_2 FILLER_166_509 ();
 sky130_fd_sc_hs__fill_2 FILLER_166_538 ();
 sky130_fd_sc_hs__fill_4 FILLER_167_0 ();
 sky130_fd_sc_hs__fill_1 FILLER_167_4 ();
 sky130_fd_sc_hs__fill_8 FILLER_167_13 ();
 sky130_fd_sc_hs__fill_8 FILLER_167_21 ();
 sky130_fd_sc_hs__fill_8 FILLER_167_29 ();
 sky130_fd_sc_hs__fill_8 FILLER_167_37 ();
 sky130_fd_sc_hs__fill_8 FILLER_167_45 ();
 sky130_fd_sc_hs__fill_4 FILLER_167_53 ();
 sky130_fd_sc_hs__fill_1 FILLER_167_57 ();
 sky130_fd_sc_hs__fill_8 FILLER_167_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_167_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_167_75 ();
 sky130_fd_sc_hs__fill_4 FILLER_167_83 ();
 sky130_fd_sc_hs__fill_1 FILLER_167_87 ();
 sky130_fd_sc_hs__fill_8 FILLER_167_94 ();
 sky130_fd_sc_hs__fill_8 FILLER_167_102 ();
 sky130_fd_sc_hs__fill_4 FILLER_167_110 ();
 sky130_fd_sc_hs__fill_2 FILLER_167_114 ();
 sky130_fd_sc_hs__fill_8 FILLER_167_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_167_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_167_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_167_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_167_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_167_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_167_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_167_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_167_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_167_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_167_213 ();
 sky130_fd_sc_hs__fill_2 FILLER_167_229 ();
 sky130_fd_sc_hs__fill_1 FILLER_167_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_167_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_167_249 ();
 sky130_fd_sc_hs__fill_4 FILLER_167_257 ();
 sky130_fd_sc_hs__fill_1 FILLER_167_261 ();
 sky130_fd_sc_hs__fill_8 FILLER_167_269 ();
 sky130_fd_sc_hs__fill_8 FILLER_167_277 ();
 sky130_fd_sc_hs__fill_4 FILLER_167_285 ();
 sky130_fd_sc_hs__fill_1 FILLER_167_289 ();
 sky130_fd_sc_hs__fill_2 FILLER_167_291 ();
 sky130_fd_sc_hs__fill_4 FILLER_167_327 ();
 sky130_fd_sc_hs__fill_2 FILLER_167_331 ();
 sky130_fd_sc_hs__fill_4 FILLER_167_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_167_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_167_357 ();
 sky130_fd_sc_hs__fill_2 FILLER_167_365 ();
 sky130_fd_sc_hs__fill_1 FILLER_167_367 ();
 sky130_fd_sc_hs__fill_2 FILLER_167_388 ();
 sky130_fd_sc_hs__fill_1 FILLER_167_390 ();
 sky130_fd_sc_hs__fill_4 FILLER_167_396 ();
 sky130_fd_sc_hs__fill_1 FILLER_167_400 ();
 sky130_fd_sc_hs__fill_1 FILLER_167_405 ();
 sky130_fd_sc_hs__fill_2 FILLER_167_413 ();
 sky130_fd_sc_hs__fill_8 FILLER_167_437 ();
 sky130_fd_sc_hs__fill_4 FILLER_167_445 ();
 sky130_fd_sc_hs__fill_2 FILLER_167_449 ();
 sky130_fd_sc_hs__fill_1 FILLER_167_451 ();
 sky130_fd_sc_hs__fill_8 FILLER_167_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_167_473 ();
 sky130_fd_sc_hs__fill_2 FILLER_167_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_167_514 ();
 sky130_fd_sc_hs__fill_8 FILLER_167_523 ();
 sky130_fd_sc_hs__fill_1 FILLER_167_531 ();
 sky130_fd_sc_hs__fill_4 FILLER_168_0 ();
 sky130_fd_sc_hs__fill_1 FILLER_168_4 ();
 sky130_fd_sc_hs__fill_8 FILLER_168_13 ();
 sky130_fd_sc_hs__fill_8 FILLER_168_21 ();
 sky130_fd_sc_hs__fill_8 FILLER_168_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_168_38 ();
 sky130_fd_sc_hs__fill_4 FILLER_168_46 ();
 sky130_fd_sc_hs__fill_2 FILLER_168_50 ();
 sky130_fd_sc_hs__fill_1 FILLER_168_52 ();
 sky130_fd_sc_hs__fill_8 FILLER_168_60 ();
 sky130_fd_sc_hs__fill_8 FILLER_168_68 ();
 sky130_fd_sc_hs__fill_8 FILLER_168_76 ();
 sky130_fd_sc_hs__fill_2 FILLER_168_84 ();
 sky130_fd_sc_hs__fill_1 FILLER_168_86 ();
 sky130_fd_sc_hs__fill_4 FILLER_168_98 ();
 sky130_fd_sc_hs__fill_2 FILLER_168_102 ();
 sky130_fd_sc_hs__fill_1 FILLER_168_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_168_111 ();
 sky130_fd_sc_hs__fill_8 FILLER_168_119 ();
 sky130_fd_sc_hs__fill_8 FILLER_168_127 ();
 sky130_fd_sc_hs__fill_8 FILLER_168_135 ();
 sky130_fd_sc_hs__fill_2 FILLER_168_143 ();
 sky130_fd_sc_hs__fill_8 FILLER_168_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_168_154 ();
 sky130_fd_sc_hs__fill_2 FILLER_168_162 ();
 sky130_fd_sc_hs__fill_1 FILLER_168_202 ();
 sky130_fd_sc_hs__fill_1 FILLER_168_224 ();
 sky130_fd_sc_hs__fill_8 FILLER_168_238 ();
 sky130_fd_sc_hs__fill_2 FILLER_168_246 ();
 sky130_fd_sc_hs__fill_1 FILLER_168_248 ();
 sky130_fd_sc_hs__fill_8 FILLER_168_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_168_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_168_278 ();
 sky130_fd_sc_hs__fill_4 FILLER_168_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_168_306 ();
 sky130_fd_sc_hs__fill_4 FILLER_168_314 ();
 sky130_fd_sc_hs__fill_1 FILLER_168_318 ();
 sky130_fd_sc_hs__fill_4 FILLER_168_320 ();
 sky130_fd_sc_hs__fill_1 FILLER_168_324 ();
 sky130_fd_sc_hs__fill_1 FILLER_168_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_168_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_168_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_168_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_168_423 ();
 sky130_fd_sc_hs__fill_4 FILLER_168_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_168_436 ();
 sky130_fd_sc_hs__fill_4 FILLER_168_444 ();
 sky130_fd_sc_hs__fill_2 FILLER_168_448 ();
 sky130_fd_sc_hs__fill_1 FILLER_168_450 ();
 sky130_fd_sc_hs__fill_8 FILLER_168_469 ();
 sky130_fd_sc_hs__fill_4 FILLER_168_477 ();
 sky130_fd_sc_hs__fill_2 FILLER_168_481 ();
 sky130_fd_sc_hs__fill_1 FILLER_168_483 ();
 sky130_fd_sc_hs__fill_4 FILLER_168_494 ();
 sky130_fd_sc_hs__fill_2 FILLER_168_498 ();
 sky130_fd_sc_hs__fill_1 FILLER_168_500 ();
 sky130_fd_sc_hs__fill_8 FILLER_168_529 ();
 sky130_fd_sc_hs__fill_2 FILLER_168_537 ();
 sky130_fd_sc_hs__fill_1 FILLER_168_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_169_0 ();
 sky130_fd_sc_hs__fill_4 FILLER_169_8 ();
 sky130_fd_sc_hs__fill_1 FILLER_169_12 ();
 sky130_fd_sc_hs__fill_8 FILLER_169_21 ();
 sky130_fd_sc_hs__fill_8 FILLER_169_29 ();
 sky130_fd_sc_hs__fill_8 FILLER_169_37 ();
 sky130_fd_sc_hs__fill_8 FILLER_169_45 ();
 sky130_fd_sc_hs__fill_4 FILLER_169_53 ();
 sky130_fd_sc_hs__fill_1 FILLER_169_57 ();
 sky130_fd_sc_hs__fill_4 FILLER_169_59 ();
 sky130_fd_sc_hs__fill_1 FILLER_169_63 ();
 sky130_fd_sc_hs__fill_2 FILLER_169_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_169_82 ();
 sky130_fd_sc_hs__fill_4 FILLER_169_100 ();
 sky130_fd_sc_hs__fill_1 FILLER_169_104 ();
 sky130_fd_sc_hs__fill_1 FILLER_169_115 ();
 sky130_fd_sc_hs__fill_1 FILLER_169_127 ();
 sky130_fd_sc_hs__fill_8 FILLER_169_131 ();
 sky130_fd_sc_hs__fill_8 FILLER_169_139 ();
 sky130_fd_sc_hs__fill_8 FILLER_169_147 ();
 sky130_fd_sc_hs__fill_8 FILLER_169_155 ();
 sky130_fd_sc_hs__fill_8 FILLER_169_163 ();
 sky130_fd_sc_hs__fill_2 FILLER_169_171 ();
 sky130_fd_sc_hs__fill_1 FILLER_169_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_169_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_169_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_169_191 ();
 sky130_fd_sc_hs__fill_2 FILLER_169_199 ();
 sky130_fd_sc_hs__fill_1 FILLER_169_201 ();
 sky130_fd_sc_hs__fill_8 FILLER_169_217 ();
 sky130_fd_sc_hs__fill_4 FILLER_169_225 ();
 sky130_fd_sc_hs__fill_2 FILLER_169_229 ();
 sky130_fd_sc_hs__fill_1 FILLER_169_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_169_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_169_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_169_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_169_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_169_265 ();
 sky130_fd_sc_hs__fill_4 FILLER_169_291 ();
 sky130_fd_sc_hs__fill_2 FILLER_169_295 ();
 sky130_fd_sc_hs__fill_1 FILLER_169_297 ();
 sky130_fd_sc_hs__fill_8 FILLER_169_309 ();
 sky130_fd_sc_hs__fill_8 FILLER_169_317 ();
 sky130_fd_sc_hs__fill_8 FILLER_169_325 ();
 sky130_fd_sc_hs__fill_2 FILLER_169_333 ();
 sky130_fd_sc_hs__fill_1 FILLER_169_335 ();
 sky130_fd_sc_hs__fill_4 FILLER_169_341 ();
 sky130_fd_sc_hs__fill_2 FILLER_169_345 ();
 sky130_fd_sc_hs__fill_1 FILLER_169_347 ();
 sky130_fd_sc_hs__fill_1 FILLER_169_349 ();
 sky130_fd_sc_hs__fill_4 FILLER_169_353 ();
 sky130_fd_sc_hs__fill_8 FILLER_169_361 ();
 sky130_fd_sc_hs__fill_8 FILLER_169_369 ();
 sky130_fd_sc_hs__fill_8 FILLER_169_377 ();
 sky130_fd_sc_hs__fill_4 FILLER_169_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_169_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_169_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_169_426 ();
 sky130_fd_sc_hs__fill_8 FILLER_169_434 ();
 sky130_fd_sc_hs__fill_4 FILLER_169_442 ();
 sky130_fd_sc_hs__fill_2 FILLER_169_446 ();
 sky130_fd_sc_hs__fill_1 FILLER_169_448 ();
 sky130_fd_sc_hs__fill_4 FILLER_169_452 ();
 sky130_fd_sc_hs__fill_1 FILLER_169_456 ();
 sky130_fd_sc_hs__fill_2 FILLER_169_461 ();
 sky130_fd_sc_hs__fill_1 FILLER_169_463 ();
 sky130_fd_sc_hs__fill_4 FILLER_169_465 ();
 sky130_fd_sc_hs__fill_2 FILLER_169_469 ();
 sky130_fd_sc_hs__fill_2 FILLER_169_479 ();
 sky130_fd_sc_hs__fill_2 FILLER_169_498 ();
 sky130_fd_sc_hs__fill_1 FILLER_169_508 ();
 sky130_fd_sc_hs__fill_4 FILLER_169_516 ();
 sky130_fd_sc_hs__fill_2 FILLER_169_520 ();
 sky130_fd_sc_hs__fill_8 FILLER_169_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_169_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_169_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_170_0 ();
 sky130_fd_sc_hs__fill_1 FILLER_170_8 ();
 sky130_fd_sc_hs__fill_4 FILLER_170_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_170_51 ();
 sky130_fd_sc_hs__fill_4 FILLER_170_59 ();
 sky130_fd_sc_hs__fill_1 FILLER_170_63 ();
 sky130_fd_sc_hs__fill_4 FILLER_170_81 ();
 sky130_fd_sc_hs__fill_2 FILLER_170_85 ();
 sky130_fd_sc_hs__fill_1 FILLER_170_88 ();
 sky130_fd_sc_hs__fill_2 FILLER_170_94 ();
 sky130_fd_sc_hs__fill_2 FILLER_170_103 ();
 sky130_fd_sc_hs__fill_2 FILLER_170_110 ();
 sky130_fd_sc_hs__fill_2 FILLER_170_119 ();
 sky130_fd_sc_hs__fill_1 FILLER_170_121 ();
 sky130_fd_sc_hs__fill_8 FILLER_170_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_170_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_170_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_170_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_170_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_170_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_170_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_170_202 ();
 sky130_fd_sc_hs__fill_1 FILLER_170_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_170_208 ();
 sky130_fd_sc_hs__fill_8 FILLER_170_216 ();
 sky130_fd_sc_hs__fill_8 FILLER_170_224 ();
 sky130_fd_sc_hs__fill_8 FILLER_170_232 ();
 sky130_fd_sc_hs__fill_8 FILLER_170_240 ();
 sky130_fd_sc_hs__fill_8 FILLER_170_248 ();
 sky130_fd_sc_hs__fill_4 FILLER_170_256 ();
 sky130_fd_sc_hs__fill_1 FILLER_170_260 ();
 sky130_fd_sc_hs__fill_4 FILLER_170_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_170_269 ();
 sky130_fd_sc_hs__fill_8 FILLER_170_277 ();
 sky130_fd_sc_hs__fill_4 FILLER_170_285 ();
 sky130_fd_sc_hs__fill_4 FILLER_170_301 ();
 sky130_fd_sc_hs__fill_8 FILLER_170_309 ();
 sky130_fd_sc_hs__fill_2 FILLER_170_317 ();
 sky130_fd_sc_hs__fill_4 FILLER_170_320 ();
 sky130_fd_sc_hs__fill_2 FILLER_170_324 ();
 sky130_fd_sc_hs__fill_8 FILLER_170_329 ();
 sky130_fd_sc_hs__fill_8 FILLER_170_337 ();
 sky130_fd_sc_hs__fill_8 FILLER_170_345 ();
 sky130_fd_sc_hs__fill_8 FILLER_170_353 ();
 sky130_fd_sc_hs__fill_4 FILLER_170_361 ();
 sky130_fd_sc_hs__fill_8 FILLER_170_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_170_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_170_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_170_386 ();
 sky130_fd_sc_hs__fill_4 FILLER_170_394 ();
 sky130_fd_sc_hs__fill_2 FILLER_170_398 ();
 sky130_fd_sc_hs__fill_1 FILLER_170_400 ();
 sky130_fd_sc_hs__fill_8 FILLER_170_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_170_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_170_434 ();
 sky130_fd_sc_hs__fill_4 FILLER_170_436 ();
 sky130_fd_sc_hs__fill_2 FILLER_170_440 ();
 sky130_fd_sc_hs__fill_1 FILLER_170_442 ();
 sky130_fd_sc_hs__fill_2 FILLER_170_467 ();
 sky130_fd_sc_hs__fill_1 FILLER_170_469 ();
 sky130_fd_sc_hs__fill_2 FILLER_170_490 ();
 sky130_fd_sc_hs__fill_1 FILLER_170_492 ();
 sky130_fd_sc_hs__fill_1 FILLER_170_494 ();
 sky130_fd_sc_hs__fill_4 FILLER_170_521 ();
 sky130_fd_sc_hs__fill_1 FILLER_170_525 ();
 sky130_fd_sc_hs__fill_4 FILLER_170_534 ();
 sky130_fd_sc_hs__fill_2 FILLER_170_538 ();
 sky130_fd_sc_hs__fill_8 FILLER_171_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_171_8 ();
 sky130_fd_sc_hs__fill_2 FILLER_171_16 ();
 sky130_fd_sc_hs__fill_1 FILLER_171_18 ();
 sky130_fd_sc_hs__fill_4 FILLER_171_53 ();
 sky130_fd_sc_hs__fill_1 FILLER_171_57 ();
 sky130_fd_sc_hs__fill_4 FILLER_171_59 ();
 sky130_fd_sc_hs__fill_2 FILLER_171_63 ();
 sky130_fd_sc_hs__fill_1 FILLER_171_65 ();
 sky130_fd_sc_hs__fill_8 FILLER_171_71 ();
 sky130_fd_sc_hs__fill_4 FILLER_171_79 ();
 sky130_fd_sc_hs__fill_1 FILLER_171_83 ();
 sky130_fd_sc_hs__fill_4 FILLER_171_130 ();
 sky130_fd_sc_hs__fill_2 FILLER_171_134 ();
 sky130_fd_sc_hs__fill_4 FILLER_171_143 ();
 sky130_fd_sc_hs__fill_2 FILLER_171_147 ();
 sky130_fd_sc_hs__fill_1 FILLER_171_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_171_163 ();
 sky130_fd_sc_hs__fill_2 FILLER_171_171 ();
 sky130_fd_sc_hs__fill_1 FILLER_171_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_171_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_171_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_171_191 ();
 sky130_fd_sc_hs__fill_4 FILLER_171_199 ();
 sky130_fd_sc_hs__fill_4 FILLER_171_226 ();
 sky130_fd_sc_hs__fill_2 FILLER_171_230 ();
 sky130_fd_sc_hs__fill_8 FILLER_171_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_171_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_171_249 ();
 sky130_fd_sc_hs__fill_4 FILLER_171_257 ();
 sky130_fd_sc_hs__fill_2 FILLER_171_261 ();
 sky130_fd_sc_hs__fill_4 FILLER_171_271 ();
 sky130_fd_sc_hs__fill_2 FILLER_171_275 ();
 sky130_fd_sc_hs__fill_2 FILLER_171_315 ();
 sky130_fd_sc_hs__fill_1 FILLER_171_317 ();
 sky130_fd_sc_hs__fill_8 FILLER_171_335 ();
 sky130_fd_sc_hs__fill_4 FILLER_171_343 ();
 sky130_fd_sc_hs__fill_1 FILLER_171_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_171_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_171_357 ();
 sky130_fd_sc_hs__fill_4 FILLER_171_365 ();
 sky130_fd_sc_hs__fill_2 FILLER_171_369 ();
 sky130_fd_sc_hs__fill_8 FILLER_171_377 ();
 sky130_fd_sc_hs__fill_8 FILLER_171_385 ();
 sky130_fd_sc_hs__fill_8 FILLER_171_393 ();
 sky130_fd_sc_hs__fill_4 FILLER_171_401 ();
 sky130_fd_sc_hs__fill_1 FILLER_171_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_171_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_171_415 ();
 sky130_fd_sc_hs__fill_1 FILLER_171_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_171_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_171_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_171_463 ();
 sky130_fd_sc_hs__fill_4 FILLER_171_465 ();
 sky130_fd_sc_hs__fill_1 FILLER_171_469 ();
 sky130_fd_sc_hs__fill_8 FILLER_171_477 ();
 sky130_fd_sc_hs__fill_2 FILLER_171_485 ();
 sky130_fd_sc_hs__fill_1 FILLER_171_487 ();
 sky130_fd_sc_hs__fill_4 FILLER_171_517 ();
 sky130_fd_sc_hs__fill_1 FILLER_171_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_171_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_171_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_171_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_172_0 ();
 sky130_fd_sc_hs__fill_1 FILLER_172_8 ();
 sky130_fd_sc_hs__fill_4 FILLER_172_25 ();
 sky130_fd_sc_hs__fill_4 FILLER_172_30 ();
 sky130_fd_sc_hs__fill_2 FILLER_172_34 ();
 sky130_fd_sc_hs__fill_1 FILLER_172_36 ();
 sky130_fd_sc_hs__fill_8 FILLER_172_42 ();
 sky130_fd_sc_hs__fill_4 FILLER_172_50 ();
 sky130_fd_sc_hs__fill_2 FILLER_172_54 ();
 sky130_fd_sc_hs__fill_4 FILLER_172_67 ();
 sky130_fd_sc_hs__fill_2 FILLER_172_84 ();
 sky130_fd_sc_hs__fill_1 FILLER_172_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_172_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_172_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_172_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_172_112 ();
 sky130_fd_sc_hs__fill_4 FILLER_172_120 ();
 sky130_fd_sc_hs__fill_2 FILLER_172_124 ();
 sky130_fd_sc_hs__fill_1 FILLER_172_126 ();
 sky130_fd_sc_hs__fill_4 FILLER_172_140 ();
 sky130_fd_sc_hs__fill_1 FILLER_172_144 ();
 sky130_fd_sc_hs__fill_4 FILLER_172_146 ();
 sky130_fd_sc_hs__fill_1 FILLER_172_150 ();
 sky130_fd_sc_hs__fill_1 FILLER_172_164 ();
 sky130_fd_sc_hs__fill_8 FILLER_172_172 ();
 sky130_fd_sc_hs__fill_8 FILLER_172_180 ();
 sky130_fd_sc_hs__fill_8 FILLER_172_188 ();
 sky130_fd_sc_hs__fill_4 FILLER_172_196 ();
 sky130_fd_sc_hs__fill_8 FILLER_172_221 ();
 sky130_fd_sc_hs__fill_8 FILLER_172_229 ();
 sky130_fd_sc_hs__fill_8 FILLER_172_237 ();
 sky130_fd_sc_hs__fill_4 FILLER_172_245 ();
 sky130_fd_sc_hs__fill_2 FILLER_172_249 ();
 sky130_fd_sc_hs__fill_1 FILLER_172_251 ();
 sky130_fd_sc_hs__fill_8 FILLER_172_262 ();
 sky130_fd_sc_hs__fill_1 FILLER_172_270 ();
 sky130_fd_sc_hs__fill_4 FILLER_172_301 ();
 sky130_fd_sc_hs__fill_1 FILLER_172_305 ();
 sky130_fd_sc_hs__fill_8 FILLER_172_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_172_328 ();
 sky130_fd_sc_hs__fill_1 FILLER_172_336 ();
 sky130_fd_sc_hs__fill_4 FILLER_172_357 ();
 sky130_fd_sc_hs__fill_2 FILLER_172_361 ();
 sky130_fd_sc_hs__fill_1 FILLER_172_363 ();
 sky130_fd_sc_hs__fill_8 FILLER_172_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_172_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_172_383 ();
 sky130_fd_sc_hs__fill_8 FILLER_172_391 ();
 sky130_fd_sc_hs__fill_8 FILLER_172_399 ();
 sky130_fd_sc_hs__fill_8 FILLER_172_407 ();
 sky130_fd_sc_hs__fill_4 FILLER_172_415 ();
 sky130_fd_sc_hs__fill_2 FILLER_172_419 ();
 sky130_fd_sc_hs__fill_1 FILLER_172_421 ();
 sky130_fd_sc_hs__fill_8 FILLER_172_427 ();
 sky130_fd_sc_hs__fill_8 FILLER_172_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_172_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_172_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_172_460 ();
 sky130_fd_sc_hs__fill_2 FILLER_172_468 ();
 sky130_fd_sc_hs__fill_4 FILLER_172_488 ();
 sky130_fd_sc_hs__fill_1 FILLER_172_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_172_517 ();
 sky130_fd_sc_hs__fill_1 FILLER_172_525 ();
 sky130_fd_sc_hs__fill_4 FILLER_172_534 ();
 sky130_fd_sc_hs__fill_2 FILLER_172_538 ();
 sky130_fd_sc_hs__fill_8 FILLER_173_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_173_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_173_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_173_24 ();
 sky130_fd_sc_hs__fill_2 FILLER_173_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_173_44 ();
 sky130_fd_sc_hs__fill_4 FILLER_173_52 ();
 sky130_fd_sc_hs__fill_2 FILLER_173_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_173_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_173_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_173_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_173_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_173_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_173_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_173_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_173_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_173_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_173_125 ();
 sky130_fd_sc_hs__fill_4 FILLER_173_133 ();
 sky130_fd_sc_hs__fill_2 FILLER_173_153 ();
 sky130_fd_sc_hs__fill_1 FILLER_173_155 ();
 sky130_fd_sc_hs__fill_8 FILLER_173_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_173_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_173_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_173_199 ();
 sky130_fd_sc_hs__fill_2 FILLER_173_207 ();
 sky130_fd_sc_hs__fill_2 FILLER_173_229 ();
 sky130_fd_sc_hs__fill_1 FILLER_173_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_173_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_173_241 ();
 sky130_fd_sc_hs__fill_2 FILLER_173_249 ();
 sky130_fd_sc_hs__fill_1 FILLER_173_251 ();
 sky130_fd_sc_hs__fill_8 FILLER_173_282 ();
 sky130_fd_sc_hs__fill_8 FILLER_173_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_173_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_173_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_173_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_173_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_173_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_173_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_173_347 ();
 sky130_fd_sc_hs__fill_4 FILLER_173_360 ();
 sky130_fd_sc_hs__fill_1 FILLER_173_364 ();
 sky130_fd_sc_hs__fill_1 FILLER_173_370 ();
 sky130_fd_sc_hs__fill_8 FILLER_173_380 ();
 sky130_fd_sc_hs__fill_8 FILLER_173_388 ();
 sky130_fd_sc_hs__fill_8 FILLER_173_396 ();
 sky130_fd_sc_hs__fill_2 FILLER_173_404 ();
 sky130_fd_sc_hs__fill_4 FILLER_173_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_173_414 ();
 sky130_fd_sc_hs__fill_2 FILLER_173_422 ();
 sky130_fd_sc_hs__fill_8 FILLER_173_429 ();
 sky130_fd_sc_hs__fill_2 FILLER_173_455 ();
 sky130_fd_sc_hs__fill_8 FILLER_173_465 ();
 sky130_fd_sc_hs__fill_1 FILLER_173_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_173_504 ();
 sky130_fd_sc_hs__fill_8 FILLER_173_512 ();
 sky130_fd_sc_hs__fill_2 FILLER_173_520 ();
 sky130_fd_sc_hs__fill_8 FILLER_173_523 ();
 sky130_fd_sc_hs__fill_1 FILLER_173_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_174_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_174_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_174_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_174_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_174_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_174_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_174_38 ();
 sky130_fd_sc_hs__fill_4 FILLER_174_46 ();
 sky130_fd_sc_hs__fill_1 FILLER_174_50 ();
 sky130_fd_sc_hs__fill_8 FILLER_174_73 ();
 sky130_fd_sc_hs__fill_4 FILLER_174_81 ();
 sky130_fd_sc_hs__fill_2 FILLER_174_85 ();
 sky130_fd_sc_hs__fill_8 FILLER_174_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_174_96 ();
 sky130_fd_sc_hs__fill_1 FILLER_174_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_174_118 ();
 sky130_fd_sc_hs__fill_8 FILLER_174_126 ();
 sky130_fd_sc_hs__fill_8 FILLER_174_134 ();
 sky130_fd_sc_hs__fill_2 FILLER_174_142 ();
 sky130_fd_sc_hs__fill_1 FILLER_174_144 ();
 sky130_fd_sc_hs__fill_4 FILLER_174_163 ();
 sky130_fd_sc_hs__fill_2 FILLER_174_167 ();
 sky130_fd_sc_hs__fill_1 FILLER_174_169 ();
 sky130_fd_sc_hs__fill_8 FILLER_174_193 ();
 sky130_fd_sc_hs__fill_2 FILLER_174_201 ();
 sky130_fd_sc_hs__fill_4 FILLER_174_204 ();
 sky130_fd_sc_hs__fill_2 FILLER_174_208 ();
 sky130_fd_sc_hs__fill_1 FILLER_174_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_174_237 ();
 sky130_fd_sc_hs__fill_8 FILLER_174_245 ();
 sky130_fd_sc_hs__fill_1 FILLER_174_253 ();
 sky130_fd_sc_hs__fill_8 FILLER_174_262 ();
 sky130_fd_sc_hs__fill_4 FILLER_174_270 ();
 sky130_fd_sc_hs__fill_4 FILLER_174_286 ();
 sky130_fd_sc_hs__fill_2 FILLER_174_290 ();
 sky130_fd_sc_hs__fill_8 FILLER_174_300 ();
 sky130_fd_sc_hs__fill_2 FILLER_174_308 ();
 sky130_fd_sc_hs__fill_1 FILLER_174_310 ();
 sky130_fd_sc_hs__fill_8 FILLER_174_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_174_328 ();
 sky130_fd_sc_hs__fill_2 FILLER_174_336 ();
 sky130_fd_sc_hs__fill_1 FILLER_174_338 ();
 sky130_fd_sc_hs__fill_8 FILLER_174_357 ();
 sky130_fd_sc_hs__fill_1 FILLER_174_365 ();
 sky130_fd_sc_hs__fill_2 FILLER_174_370 ();
 sky130_fd_sc_hs__fill_2 FILLER_174_384 ();
 sky130_fd_sc_hs__fill_4 FILLER_174_397 ();
 sky130_fd_sc_hs__fill_2 FILLER_174_401 ();
 sky130_fd_sc_hs__fill_1 FILLER_174_403 ();
 sky130_fd_sc_hs__fill_8 FILLER_174_419 ();
 sky130_fd_sc_hs__fill_8 FILLER_174_427 ();
 sky130_fd_sc_hs__fill_8 FILLER_174_436 ();
 sky130_fd_sc_hs__fill_1 FILLER_174_444 ();
 sky130_fd_sc_hs__fill_2 FILLER_174_490 ();
 sky130_fd_sc_hs__fill_1 FILLER_174_492 ();
 sky130_fd_sc_hs__fill_4 FILLER_174_498 ();
 sky130_fd_sc_hs__fill_8 FILLER_175_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_175_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_175_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_175_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_175_37 ();
 sky130_fd_sc_hs__fill_2 FILLER_175_45 ();
 sky130_fd_sc_hs__fill_1 FILLER_175_47 ();
 sky130_fd_sc_hs__fill_8 FILLER_175_72 ();
 sky130_fd_sc_hs__fill_2 FILLER_175_80 ();
 sky130_fd_sc_hs__fill_1 FILLER_175_98 ();
 sky130_fd_sc_hs__fill_2 FILLER_175_114 ();
 sky130_fd_sc_hs__fill_2 FILLER_175_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_175_122 ();
 sky130_fd_sc_hs__fill_8 FILLER_175_130 ();
 sky130_fd_sc_hs__fill_4 FILLER_175_138 ();
 sky130_fd_sc_hs__fill_2 FILLER_175_142 ();
 sky130_fd_sc_hs__fill_1 FILLER_175_144 ();
 sky130_fd_sc_hs__fill_1 FILLER_175_150 ();
 sky130_fd_sc_hs__fill_8 FILLER_175_164 ();
 sky130_fd_sc_hs__fill_2 FILLER_175_172 ();
 sky130_fd_sc_hs__fill_2 FILLER_175_189 ();
 sky130_fd_sc_hs__fill_8 FILLER_175_195 ();
 sky130_fd_sc_hs__fill_8 FILLER_175_203 ();
 sky130_fd_sc_hs__fill_8 FILLER_175_211 ();
 sky130_fd_sc_hs__fill_8 FILLER_175_219 ();
 sky130_fd_sc_hs__fill_4 FILLER_175_227 ();
 sky130_fd_sc_hs__fill_1 FILLER_175_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_175_233 ();
 sky130_fd_sc_hs__fill_4 FILLER_175_241 ();
 sky130_fd_sc_hs__fill_1 FILLER_175_245 ();
 sky130_fd_sc_hs__fill_8 FILLER_175_258 ();
 sky130_fd_sc_hs__fill_8 FILLER_175_266 ();
 sky130_fd_sc_hs__fill_8 FILLER_175_274 ();
 sky130_fd_sc_hs__fill_8 FILLER_175_282 ();
 sky130_fd_sc_hs__fill_8 FILLER_175_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_175_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_175_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_175_315 ();
 sky130_fd_sc_hs__fill_4 FILLER_175_323 ();
 sky130_fd_sc_hs__fill_4 FILLER_175_349 ();
 sky130_fd_sc_hs__fill_4 FILLER_175_362 ();
 sky130_fd_sc_hs__fill_1 FILLER_175_383 ();
 sky130_fd_sc_hs__fill_8 FILLER_175_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_175_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_175_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_175_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_175_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_175_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_175_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_175_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_175_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_175_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_175_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_175_465 ();
 sky130_fd_sc_hs__fill_1 FILLER_175_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_175_478 ();
 sky130_fd_sc_hs__fill_8 FILLER_175_486 ();
 sky130_fd_sc_hs__fill_1 FILLER_175_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_175_498 ();
 sky130_fd_sc_hs__fill_8 FILLER_175_514 ();
 sky130_fd_sc_hs__fill_8 FILLER_175_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_175_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_175_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_176_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_176_8 ();
 sky130_fd_sc_hs__fill_2 FILLER_176_16 ();
 sky130_fd_sc_hs__fill_1 FILLER_176_18 ();
 sky130_fd_sc_hs__fill_8 FILLER_176_37 ();
 sky130_fd_sc_hs__fill_8 FILLER_176_45 ();
 sky130_fd_sc_hs__fill_4 FILLER_176_53 ();
 sky130_fd_sc_hs__fill_2 FILLER_176_57 ();
 sky130_fd_sc_hs__fill_2 FILLER_176_64 ();
 sky130_fd_sc_hs__fill_1 FILLER_176_66 ();
 sky130_fd_sc_hs__fill_8 FILLER_176_74 ();
 sky130_fd_sc_hs__fill_4 FILLER_176_82 ();
 sky130_fd_sc_hs__fill_1 FILLER_176_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_176_103 ();
 sky130_fd_sc_hs__fill_8 FILLER_176_131 ();
 sky130_fd_sc_hs__fill_4 FILLER_176_139 ();
 sky130_fd_sc_hs__fill_2 FILLER_176_143 ();
 sky130_fd_sc_hs__fill_8 FILLER_176_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_176_154 ();
 sky130_fd_sc_hs__fill_4 FILLER_176_162 ();
 sky130_fd_sc_hs__fill_2 FILLER_176_166 ();
 sky130_fd_sc_hs__fill_1 FILLER_176_168 ();
 sky130_fd_sc_hs__fill_2 FILLER_176_201 ();
 sky130_fd_sc_hs__fill_8 FILLER_176_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_176_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_176_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_176_228 ();
 sky130_fd_sc_hs__fill_2 FILLER_176_236 ();
 sky130_fd_sc_hs__fill_1 FILLER_176_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_176_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_176_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_176_278 ();
 sky130_fd_sc_hs__fill_2 FILLER_176_286 ();
 sky130_fd_sc_hs__fill_1 FILLER_176_288 ();
 sky130_fd_sc_hs__fill_8 FILLER_176_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_176_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_176_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_176_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_176_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_176_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_176_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_176_376 ();
 sky130_fd_sc_hs__fill_2 FILLER_176_378 ();
 sky130_fd_sc_hs__fill_4 FILLER_176_401 ();
 sky130_fd_sc_hs__fill_2 FILLER_176_405 ();
 sky130_fd_sc_hs__fill_1 FILLER_176_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_176_420 ();
 sky130_fd_sc_hs__fill_4 FILLER_176_428 ();
 sky130_fd_sc_hs__fill_2 FILLER_176_432 ();
 sky130_fd_sc_hs__fill_1 FILLER_176_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_176_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_176_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_176_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_176_460 ();
 sky130_fd_sc_hs__fill_4 FILLER_176_468 ();
 sky130_fd_sc_hs__fill_1 FILLER_176_472 ();
 sky130_fd_sc_hs__fill_8 FILLER_176_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_176_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_176_492 ();
 sky130_fd_sc_hs__fill_4 FILLER_176_517 ();
 sky130_fd_sc_hs__fill_2 FILLER_176_521 ();
 sky130_fd_sc_hs__fill_1 FILLER_176_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_176_532 ();
 sky130_fd_sc_hs__fill_8 FILLER_177_0 ();
 sky130_fd_sc_hs__fill_4 FILLER_177_8 ();
 sky130_fd_sc_hs__fill_1 FILLER_177_12 ();
 sky130_fd_sc_hs__fill_4 FILLER_177_21 ();
 sky130_fd_sc_hs__fill_8 FILLER_177_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_177_46 ();
 sky130_fd_sc_hs__fill_4 FILLER_177_54 ();
 sky130_fd_sc_hs__fill_4 FILLER_177_59 ();
 sky130_fd_sc_hs__fill_2 FILLER_177_63 ();
 sky130_fd_sc_hs__fill_8 FILLER_177_78 ();
 sky130_fd_sc_hs__fill_4 FILLER_177_86 ();
 sky130_fd_sc_hs__fill_1 FILLER_177_90 ();
 sky130_fd_sc_hs__fill_1 FILLER_177_98 ();
 sky130_fd_sc_hs__fill_8 FILLER_177_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_177_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_177_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_177_125 ();
 sky130_fd_sc_hs__fill_2 FILLER_177_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_177_158 ();
 sky130_fd_sc_hs__fill_8 FILLER_177_166 ();
 sky130_fd_sc_hs__fill_8 FILLER_177_175 ();
 sky130_fd_sc_hs__fill_1 FILLER_177_183 ();
 sky130_fd_sc_hs__fill_2 FILLER_177_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_177_206 ();
 sky130_fd_sc_hs__fill_8 FILLER_177_214 ();
 sky130_fd_sc_hs__fill_8 FILLER_177_222 ();
 sky130_fd_sc_hs__fill_2 FILLER_177_230 ();
 sky130_fd_sc_hs__fill_8 FILLER_177_233 ();
 sky130_fd_sc_hs__fill_4 FILLER_177_241 ();
 sky130_fd_sc_hs__fill_2 FILLER_177_245 ();
 sky130_fd_sc_hs__fill_8 FILLER_177_277 ();
 sky130_fd_sc_hs__fill_4 FILLER_177_285 ();
 sky130_fd_sc_hs__fill_1 FILLER_177_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_177_325 ();
 sky130_fd_sc_hs__fill_8 FILLER_177_333 ();
 sky130_fd_sc_hs__fill_4 FILLER_177_341 ();
 sky130_fd_sc_hs__fill_2 FILLER_177_345 ();
 sky130_fd_sc_hs__fill_1 FILLER_177_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_177_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_177_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_177_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_177_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_177_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_177_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_177_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_177_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_177_407 ();
 sky130_fd_sc_hs__fill_2 FILLER_177_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_177_422 ();
 sky130_fd_sc_hs__fill_2 FILLER_177_430 ();
 sky130_fd_sc_hs__fill_1 FILLER_177_432 ();
 sky130_fd_sc_hs__fill_8 FILLER_177_445 ();
 sky130_fd_sc_hs__fill_8 FILLER_177_453 ();
 sky130_fd_sc_hs__fill_2 FILLER_177_461 ();
 sky130_fd_sc_hs__fill_1 FILLER_177_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_177_488 ();
 sky130_fd_sc_hs__fill_2 FILLER_177_496 ();
 sky130_fd_sc_hs__fill_8 FILLER_177_506 ();
 sky130_fd_sc_hs__fill_8 FILLER_177_514 ();
 sky130_fd_sc_hs__fill_8 FILLER_177_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_177_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_177_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_178_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_178_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_178_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_178_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_178_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_178_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_178_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_178_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_178_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_178_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_178_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_178_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_178_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_178_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_178_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_178_104 ();
 sky130_fd_sc_hs__fill_4 FILLER_178_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_178_132 ();
 sky130_fd_sc_hs__fill_4 FILLER_178_140 ();
 sky130_fd_sc_hs__fill_1 FILLER_178_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_178_156 ();
 sky130_fd_sc_hs__fill_8 FILLER_178_164 ();
 sky130_fd_sc_hs__fill_8 FILLER_178_172 ();
 sky130_fd_sc_hs__fill_8 FILLER_178_180 ();
 sky130_fd_sc_hs__fill_8 FILLER_178_188 ();
 sky130_fd_sc_hs__fill_4 FILLER_178_196 ();
 sky130_fd_sc_hs__fill_2 FILLER_178_200 ();
 sky130_fd_sc_hs__fill_1 FILLER_178_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_178_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_178_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_178_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_178_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_178_236 ();
 sky130_fd_sc_hs__fill_4 FILLER_178_244 ();
 sky130_fd_sc_hs__fill_1 FILLER_178_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_178_270 ();
 sky130_fd_sc_hs__fill_2 FILLER_178_278 ();
 sky130_fd_sc_hs__fill_1 FILLER_178_280 ();
 sky130_fd_sc_hs__fill_8 FILLER_178_290 ();
 sky130_fd_sc_hs__fill_8 FILLER_178_298 ();
 sky130_fd_sc_hs__fill_8 FILLER_178_306 ();
 sky130_fd_sc_hs__fill_4 FILLER_178_314 ();
 sky130_fd_sc_hs__fill_1 FILLER_178_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_178_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_178_328 ();
 sky130_fd_sc_hs__fill_2 FILLER_178_336 ();
 sky130_fd_sc_hs__fill_1 FILLER_178_338 ();
 sky130_fd_sc_hs__fill_8 FILLER_178_366 ();
 sky130_fd_sc_hs__fill_2 FILLER_178_374 ();
 sky130_fd_sc_hs__fill_1 FILLER_178_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_178_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_178_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_178_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_178_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_178_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_178_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_178_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_178_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_178_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_178_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_178_452 ();
 sky130_fd_sc_hs__fill_2 FILLER_178_460 ();
 sky130_fd_sc_hs__fill_1 FILLER_178_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_178_494 ();
 sky130_fd_sc_hs__fill_2 FILLER_178_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_178_516 ();
 sky130_fd_sc_hs__fill_8 FILLER_178_532 ();
 sky130_fd_sc_hs__fill_8 FILLER_179_0 ();
 sky130_fd_sc_hs__fill_2 FILLER_179_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_179_18 ();
 sky130_fd_sc_hs__fill_8 FILLER_179_26 ();
 sky130_fd_sc_hs__fill_8 FILLER_179_34 ();
 sky130_fd_sc_hs__fill_8 FILLER_179_42 ();
 sky130_fd_sc_hs__fill_8 FILLER_179_50 ();
 sky130_fd_sc_hs__fill_8 FILLER_179_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_179_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_179_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_179_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_179_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_179_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_179_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_179_115 ();
 sky130_fd_sc_hs__fill_4 FILLER_179_134 ();
 sky130_fd_sc_hs__fill_2 FILLER_179_138 ();
 sky130_fd_sc_hs__fill_4 FILLER_179_145 ();
 sky130_fd_sc_hs__fill_2 FILLER_179_149 ();
 sky130_fd_sc_hs__fill_1 FILLER_179_151 ();
 sky130_fd_sc_hs__fill_8 FILLER_179_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_179_173 ();
 sky130_fd_sc_hs__fill_4 FILLER_179_175 ();
 sky130_fd_sc_hs__fill_2 FILLER_179_179 ();
 sky130_fd_sc_hs__fill_1 FILLER_179_181 ();
 sky130_fd_sc_hs__fill_8 FILLER_179_185 ();
 sky130_fd_sc_hs__fill_8 FILLER_179_193 ();
 sky130_fd_sc_hs__fill_4 FILLER_179_201 ();
 sky130_fd_sc_hs__fill_2 FILLER_179_205 ();
 sky130_fd_sc_hs__fill_1 FILLER_179_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_179_211 ();
 sky130_fd_sc_hs__fill_8 FILLER_179_219 ();
 sky130_fd_sc_hs__fill_4 FILLER_179_227 ();
 sky130_fd_sc_hs__fill_1 FILLER_179_231 ();
 sky130_fd_sc_hs__fill_4 FILLER_179_233 ();
 sky130_fd_sc_hs__fill_2 FILLER_179_237 ();
 sky130_fd_sc_hs__fill_8 FILLER_179_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_179_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_179_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_179_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_179_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_179_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_179_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_179_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_179_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_179_347 ();
 sky130_fd_sc_hs__fill_2 FILLER_179_367 ();
 sky130_fd_sc_hs__fill_1 FILLER_179_369 ();
 sky130_fd_sc_hs__fill_8 FILLER_179_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_179_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_179_394 ();
 sky130_fd_sc_hs__fill_4 FILLER_179_402 ();
 sky130_fd_sc_hs__fill_2 FILLER_179_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_179_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_179_426 ();
 sky130_fd_sc_hs__fill_8 FILLER_179_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_179_442 ();
 sky130_fd_sc_hs__fill_8 FILLER_179_450 ();
 sky130_fd_sc_hs__fill_4 FILLER_179_458 ();
 sky130_fd_sc_hs__fill_2 FILLER_179_462 ();
 sky130_fd_sc_hs__fill_8 FILLER_179_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_179_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_179_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_179_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_179_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_179_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_179_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_179_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_179_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_179_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_179_539 ();
 sky130_fd_sc_hs__fill_4 FILLER_180_0 ();
 sky130_fd_sc_hs__fill_1 FILLER_180_4 ();
 sky130_fd_sc_hs__fill_8 FILLER_180_13 ();
 sky130_fd_sc_hs__fill_8 FILLER_180_21 ();
 sky130_fd_sc_hs__fill_8 FILLER_180_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_180_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_180_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_180_54 ();
 sky130_fd_sc_hs__fill_1 FILLER_180_62 ();
 sky130_fd_sc_hs__fill_4 FILLER_180_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_180_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_180_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_180_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_180_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_180_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_180_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_180_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_180_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_180_159 ();
 sky130_fd_sc_hs__fill_8 FILLER_180_167 ();
 sky130_fd_sc_hs__fill_2 FILLER_180_175 ();
 sky130_fd_sc_hs__fill_1 FILLER_180_177 ();
 sky130_fd_sc_hs__fill_1 FILLER_180_181 ();
 sky130_fd_sc_hs__fill_1 FILLER_180_204 ();
 sky130_fd_sc_hs__fill_4 FILLER_180_218 ();
 sky130_fd_sc_hs__fill_1 FILLER_180_222 ();
 sky130_fd_sc_hs__fill_8 FILLER_180_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_180_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_180_262 ();
 sky130_fd_sc_hs__fill_4 FILLER_180_270 ();
 sky130_fd_sc_hs__fill_2 FILLER_180_274 ();
 sky130_fd_sc_hs__fill_1 FILLER_180_276 ();
 sky130_fd_sc_hs__fill_8 FILLER_180_296 ();
 sky130_fd_sc_hs__fill_2 FILLER_180_304 ();
 sky130_fd_sc_hs__fill_1 FILLER_180_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_180_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_180_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_180_336 ();
 sky130_fd_sc_hs__fill_4 FILLER_180_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_180_357 ();
 sky130_fd_sc_hs__fill_4 FILLER_180_365 ();
 sky130_fd_sc_hs__fill_1 FILLER_180_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_180_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_180_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_180_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_180_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_180_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_180_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_180_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_180_434 ();
 sky130_fd_sc_hs__fill_4 FILLER_180_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_180_458 ();
 sky130_fd_sc_hs__fill_8 FILLER_180_466 ();
 sky130_fd_sc_hs__fill_8 FILLER_180_474 ();
 sky130_fd_sc_hs__fill_8 FILLER_180_482 ();
 sky130_fd_sc_hs__fill_2 FILLER_180_490 ();
 sky130_fd_sc_hs__fill_1 FILLER_180_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_180_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_180_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_180_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_180_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_180_526 ();
 sky130_fd_sc_hs__fill_4 FILLER_180_534 ();
 sky130_fd_sc_hs__fill_2 FILLER_180_538 ();
 sky130_fd_sc_hs__fill_8 FILLER_181_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_181_8 ();
 sky130_fd_sc_hs__fill_2 FILLER_181_16 ();
 sky130_fd_sc_hs__fill_2 FILLER_181_26 ();
 sky130_fd_sc_hs__fill_8 FILLER_181_47 ();
 sky130_fd_sc_hs__fill_2 FILLER_181_55 ();
 sky130_fd_sc_hs__fill_1 FILLER_181_57 ();
 sky130_fd_sc_hs__fill_1 FILLER_181_59 ();
 sky130_fd_sc_hs__fill_2 FILLER_181_65 ();
 sky130_fd_sc_hs__fill_8 FILLER_181_80 ();
 sky130_fd_sc_hs__fill_8 FILLER_181_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_181_96 ();
 sky130_fd_sc_hs__fill_4 FILLER_181_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_181_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_181_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_181_136 ();
 sky130_fd_sc_hs__fill_8 FILLER_181_144 ();
 sky130_fd_sc_hs__fill_4 FILLER_181_152 ();
 sky130_fd_sc_hs__fill_2 FILLER_181_172 ();
 sky130_fd_sc_hs__fill_4 FILLER_181_175 ();
 sky130_fd_sc_hs__fill_1 FILLER_181_179 ();
 sky130_fd_sc_hs__fill_1 FILLER_181_201 ();
 sky130_fd_sc_hs__fill_2 FILLER_181_212 ();
 sky130_fd_sc_hs__fill_1 FILLER_181_214 ();
 sky130_fd_sc_hs__fill_2 FILLER_181_230 ();
 sky130_fd_sc_hs__fill_8 FILLER_181_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_181_241 ();
 sky130_fd_sc_hs__fill_2 FILLER_181_249 ();
 sky130_fd_sc_hs__fill_1 FILLER_181_251 ();
 sky130_fd_sc_hs__fill_4 FILLER_181_255 ();
 sky130_fd_sc_hs__fill_2 FILLER_181_259 ();
 sky130_fd_sc_hs__fill_1 FILLER_181_261 ();
 sky130_fd_sc_hs__fill_8 FILLER_181_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_181_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_181_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_181_291 ();
 sky130_fd_sc_hs__fill_4 FILLER_181_332 ();
 sky130_fd_sc_hs__fill_2 FILLER_181_336 ();
 sky130_fd_sc_hs__fill_4 FILLER_181_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_181_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_181_357 ();
 sky130_fd_sc_hs__fill_4 FILLER_181_365 ();
 sky130_fd_sc_hs__fill_2 FILLER_181_369 ();
 sky130_fd_sc_hs__fill_1 FILLER_181_371 ();
 sky130_fd_sc_hs__fill_2 FILLER_181_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_181_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_181_394 ();
 sky130_fd_sc_hs__fill_4 FILLER_181_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_181_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_181_428 ();
 sky130_fd_sc_hs__fill_8 FILLER_181_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_181_444 ();
 sky130_fd_sc_hs__fill_2 FILLER_181_452 ();
 sky130_fd_sc_hs__fill_1 FILLER_181_454 ();
 sky130_fd_sc_hs__fill_1 FILLER_181_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_181_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_181_498 ();
 sky130_fd_sc_hs__fill_8 FILLER_181_506 ();
 sky130_fd_sc_hs__fill_8 FILLER_181_514 ();
 sky130_fd_sc_hs__fill_4 FILLER_181_523 ();
 sky130_fd_sc_hs__fill_1 FILLER_181_527 ();
 sky130_fd_sc_hs__fill_4 FILLER_181_536 ();
 sky130_fd_sc_hs__fill_8 FILLER_182_0 ();
 sky130_fd_sc_hs__fill_4 FILLER_182_8 ();
 sky130_fd_sc_hs__fill_1 FILLER_182_12 ();
 sky130_fd_sc_hs__fill_8 FILLER_182_21 ();
 sky130_fd_sc_hs__fill_8 FILLER_182_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_182_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_182_46 ();
 sky130_fd_sc_hs__fill_2 FILLER_182_54 ();
 sky130_fd_sc_hs__fill_1 FILLER_182_66 ();
 sky130_fd_sc_hs__fill_2 FILLER_182_84 ();
 sky130_fd_sc_hs__fill_1 FILLER_182_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_182_88 ();
 sky130_fd_sc_hs__fill_4 FILLER_182_96 ();
 sky130_fd_sc_hs__fill_2 FILLER_182_100 ();
 sky130_fd_sc_hs__fill_8 FILLER_182_122 ();
 sky130_fd_sc_hs__fill_2 FILLER_182_130 ();
 sky130_fd_sc_hs__fill_1 FILLER_182_132 ();
 sky130_fd_sc_hs__fill_4 FILLER_182_138 ();
 sky130_fd_sc_hs__fill_2 FILLER_182_142 ();
 sky130_fd_sc_hs__fill_1 FILLER_182_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_182_146 ();
 sky130_fd_sc_hs__fill_2 FILLER_182_154 ();
 sky130_fd_sc_hs__fill_4 FILLER_182_173 ();
 sky130_fd_sc_hs__fill_2 FILLER_182_177 ();
 sky130_fd_sc_hs__fill_1 FILLER_182_179 ();
 sky130_fd_sc_hs__fill_8 FILLER_182_185 ();
 sky130_fd_sc_hs__fill_8 FILLER_182_193 ();
 sky130_fd_sc_hs__fill_2 FILLER_182_201 ();
 sky130_fd_sc_hs__fill_1 FILLER_182_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_182_211 ();
 sky130_fd_sc_hs__fill_8 FILLER_182_219 ();
 sky130_fd_sc_hs__fill_8 FILLER_182_227 ();
 sky130_fd_sc_hs__fill_8 FILLER_182_235 ();
 sky130_fd_sc_hs__fill_8 FILLER_182_243 ();
 sky130_fd_sc_hs__fill_1 FILLER_182_251 ();
 sky130_fd_sc_hs__fill_4 FILLER_182_262 ();
 sky130_fd_sc_hs__fill_1 FILLER_182_266 ();
 sky130_fd_sc_hs__fill_8 FILLER_182_285 ();
 sky130_fd_sc_hs__fill_1 FILLER_182_293 ();
 sky130_fd_sc_hs__fill_2 FILLER_182_316 ();
 sky130_fd_sc_hs__fill_1 FILLER_182_318 ();
 sky130_fd_sc_hs__fill_4 FILLER_182_332 ();
 sky130_fd_sc_hs__fill_2 FILLER_182_336 ();
 sky130_fd_sc_hs__fill_4 FILLER_182_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_182_389 ();
 sky130_fd_sc_hs__fill_1 FILLER_182_400 ();
 sky130_fd_sc_hs__fill_8 FILLER_182_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_182_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_182_423 ();
 sky130_fd_sc_hs__fill_4 FILLER_182_431 ();
 sky130_fd_sc_hs__fill_2 FILLER_182_436 ();
 sky130_fd_sc_hs__fill_2 FILLER_182_459 ();
 sky130_fd_sc_hs__fill_1 FILLER_182_461 ();
 sky130_fd_sc_hs__fill_4 FILLER_182_466 ();
 sky130_fd_sc_hs__fill_1 FILLER_182_470 ();
 sky130_fd_sc_hs__fill_4 FILLER_182_498 ();
 sky130_fd_sc_hs__fill_2 FILLER_182_502 ();
 sky130_fd_sc_hs__fill_1 FILLER_182_504 ();
 sky130_fd_sc_hs__fill_8 FILLER_182_513 ();
 sky130_fd_sc_hs__fill_8 FILLER_182_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_182_529 ();
 sky130_fd_sc_hs__fill_2 FILLER_182_537 ();
 sky130_fd_sc_hs__fill_1 FILLER_182_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_183_0 ();
 sky130_fd_sc_hs__fill_4 FILLER_183_8 ();
 sky130_fd_sc_hs__fill_1 FILLER_183_12 ();
 sky130_fd_sc_hs__fill_8 FILLER_183_21 ();
 sky130_fd_sc_hs__fill_8 FILLER_183_29 ();
 sky130_fd_sc_hs__fill_8 FILLER_183_37 ();
 sky130_fd_sc_hs__fill_8 FILLER_183_45 ();
 sky130_fd_sc_hs__fill_4 FILLER_183_53 ();
 sky130_fd_sc_hs__fill_1 FILLER_183_57 ();
 sky130_fd_sc_hs__fill_8 FILLER_183_69 ();
 sky130_fd_sc_hs__fill_4 FILLER_183_77 ();
 sky130_fd_sc_hs__fill_1 FILLER_183_87 ();
 sky130_fd_sc_hs__fill_1 FILLER_183_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_183_139 ();
 sky130_fd_sc_hs__fill_8 FILLER_183_147 ();
 sky130_fd_sc_hs__fill_2 FILLER_183_155 ();
 sky130_fd_sc_hs__fill_4 FILLER_183_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_183_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_183_183 ();
 sky130_fd_sc_hs__fill_4 FILLER_183_191 ();
 sky130_fd_sc_hs__fill_1 FILLER_183_195 ();
 sky130_fd_sc_hs__fill_8 FILLER_183_201 ();
 sky130_fd_sc_hs__fill_8 FILLER_183_209 ();
 sky130_fd_sc_hs__fill_8 FILLER_183_217 ();
 sky130_fd_sc_hs__fill_4 FILLER_183_225 ();
 sky130_fd_sc_hs__fill_2 FILLER_183_229 ();
 sky130_fd_sc_hs__fill_1 FILLER_183_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_183_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_183_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_183_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_183_257 ();
 sky130_fd_sc_hs__fill_2 FILLER_183_265 ();
 sky130_fd_sc_hs__fill_1 FILLER_183_267 ();
 sky130_fd_sc_hs__fill_2 FILLER_183_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_183_283 ();
 sky130_fd_sc_hs__fill_4 FILLER_183_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_183_310 ();
 sky130_fd_sc_hs__fill_4 FILLER_183_318 ();
 sky130_fd_sc_hs__fill_1 FILLER_183_322 ();
 sky130_fd_sc_hs__fill_8 FILLER_183_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_183_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_183_347 ();
 sky130_fd_sc_hs__fill_2 FILLER_183_349 ();
 sky130_fd_sc_hs__fill_1 FILLER_183_351 ();
 sky130_fd_sc_hs__fill_4 FILLER_183_361 ();
 sky130_fd_sc_hs__fill_1 FILLER_183_365 ();
 sky130_fd_sc_hs__fill_4 FILLER_183_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_183_419 ();
 sky130_fd_sc_hs__fill_4 FILLER_183_427 ();
 sky130_fd_sc_hs__fill_2 FILLER_183_431 ();
 sky130_fd_sc_hs__fill_1 FILLER_183_433 ();
 sky130_fd_sc_hs__fill_4 FILLER_183_457 ();
 sky130_fd_sc_hs__fill_2 FILLER_183_461 ();
 sky130_fd_sc_hs__fill_1 FILLER_183_463 ();
 sky130_fd_sc_hs__fill_4 FILLER_183_465 ();
 sky130_fd_sc_hs__fill_1 FILLER_183_472 ();
 sky130_fd_sc_hs__fill_4 FILLER_183_502 ();
 sky130_fd_sc_hs__fill_1 FILLER_183_506 ();
 sky130_fd_sc_hs__fill_4 FILLER_183_515 ();
 sky130_fd_sc_hs__fill_2 FILLER_183_519 ();
 sky130_fd_sc_hs__fill_1 FILLER_183_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_183_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_183_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_183_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_184_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_184_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_184_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_184_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_184_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_184_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_184_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_184_46 ();
 sky130_fd_sc_hs__fill_4 FILLER_184_54 ();
 sky130_fd_sc_hs__fill_1 FILLER_184_58 ();
 sky130_fd_sc_hs__fill_8 FILLER_184_63 ();
 sky130_fd_sc_hs__fill_8 FILLER_184_71 ();
 sky130_fd_sc_hs__fill_8 FILLER_184_79 ();
 sky130_fd_sc_hs__fill_8 FILLER_184_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_184_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_184_104 ();
 sky130_fd_sc_hs__fill_4 FILLER_184_112 ();
 sky130_fd_sc_hs__fill_2 FILLER_184_143 ();
 sky130_fd_sc_hs__fill_8 FILLER_184_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_184_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_184_162 ();
 sky130_fd_sc_hs__fill_4 FILLER_184_170 ();
 sky130_fd_sc_hs__fill_2 FILLER_184_174 ();
 sky130_fd_sc_hs__fill_4 FILLER_184_182 ();
 sky130_fd_sc_hs__fill_1 FILLER_184_186 ();
 sky130_fd_sc_hs__fill_4 FILLER_184_190 ();
 sky130_fd_sc_hs__fill_1 FILLER_184_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_184_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_184_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_184_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_184_228 ();
 sky130_fd_sc_hs__fill_2 FILLER_184_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_184_250 ();
 sky130_fd_sc_hs__fill_2 FILLER_184_258 ();
 sky130_fd_sc_hs__fill_1 FILLER_184_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_184_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_184_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_184_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_184_286 ();
 sky130_fd_sc_hs__fill_4 FILLER_184_294 ();
 sky130_fd_sc_hs__fill_1 FILLER_184_298 ();
 sky130_fd_sc_hs__fill_8 FILLER_184_304 ();
 sky130_fd_sc_hs__fill_4 FILLER_184_312 ();
 sky130_fd_sc_hs__fill_2 FILLER_184_316 ();
 sky130_fd_sc_hs__fill_1 FILLER_184_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_184_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_184_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_184_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_184_344 ();
 sky130_fd_sc_hs__fill_2 FILLER_184_352 ();
 sky130_fd_sc_hs__fill_1 FILLER_184_354 ();
 sky130_fd_sc_hs__fill_8 FILLER_184_367 ();
 sky130_fd_sc_hs__fill_2 FILLER_184_375 ();
 sky130_fd_sc_hs__fill_8 FILLER_184_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_184_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_184_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_184_422 ();
 sky130_fd_sc_hs__fill_4 FILLER_184_430 ();
 sky130_fd_sc_hs__fill_1 FILLER_184_434 ();
 sky130_fd_sc_hs__fill_1 FILLER_184_482 ();
 sky130_fd_sc_hs__fill_4 FILLER_184_487 ();
 sky130_fd_sc_hs__fill_2 FILLER_184_491 ();
 sky130_fd_sc_hs__fill_4 FILLER_184_494 ();
 sky130_fd_sc_hs__fill_1 FILLER_184_498 ();
 sky130_fd_sc_hs__fill_8 FILLER_184_530 ();
 sky130_fd_sc_hs__fill_2 FILLER_184_538 ();
 sky130_fd_sc_hs__fill_8 FILLER_185_0 ();
 sky130_fd_sc_hs__fill_2 FILLER_185_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_185_18 ();
 sky130_fd_sc_hs__fill_8 FILLER_185_26 ();
 sky130_fd_sc_hs__fill_8 FILLER_185_34 ();
 sky130_fd_sc_hs__fill_8 FILLER_185_42 ();
 sky130_fd_sc_hs__fill_8 FILLER_185_50 ();
 sky130_fd_sc_hs__fill_4 FILLER_185_59 ();
 sky130_fd_sc_hs__fill_1 FILLER_185_63 ();
 sky130_fd_sc_hs__fill_2 FILLER_185_69 ();
 sky130_fd_sc_hs__fill_1 FILLER_185_71 ();
 sky130_fd_sc_hs__fill_4 FILLER_185_92 ();
 sky130_fd_sc_hs__fill_2 FILLER_185_96 ();
 sky130_fd_sc_hs__fill_1 FILLER_185_98 ();
 sky130_fd_sc_hs__fill_8 FILLER_185_105 ();
 sky130_fd_sc_hs__fill_2 FILLER_185_113 ();
 sky130_fd_sc_hs__fill_1 FILLER_185_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_185_117 ();
 sky130_fd_sc_hs__fill_4 FILLER_185_125 ();
 sky130_fd_sc_hs__fill_1 FILLER_185_129 ();
 sky130_fd_sc_hs__fill_8 FILLER_185_142 ();
 sky130_fd_sc_hs__fill_8 FILLER_185_156 ();
 sky130_fd_sc_hs__fill_8 FILLER_185_164 ();
 sky130_fd_sc_hs__fill_2 FILLER_185_172 ();
 sky130_fd_sc_hs__fill_4 FILLER_185_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_185_201 ();
 sky130_fd_sc_hs__fill_8 FILLER_185_209 ();
 sky130_fd_sc_hs__fill_8 FILLER_185_217 ();
 sky130_fd_sc_hs__fill_4 FILLER_185_225 ();
 sky130_fd_sc_hs__fill_2 FILLER_185_229 ();
 sky130_fd_sc_hs__fill_1 FILLER_185_231 ();
 sky130_fd_sc_hs__fill_2 FILLER_185_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_185_243 ();
 sky130_fd_sc_hs__fill_8 FILLER_185_251 ();
 sky130_fd_sc_hs__fill_2 FILLER_185_259 ();
 sky130_fd_sc_hs__fill_8 FILLER_185_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_185_273 ();
 sky130_fd_sc_hs__fill_4 FILLER_185_281 ();
 sky130_fd_sc_hs__fill_2 FILLER_185_291 ();
 sky130_fd_sc_hs__fill_1 FILLER_185_293 ();
 sky130_fd_sc_hs__fill_8 FILLER_185_302 ();
 sky130_fd_sc_hs__fill_8 FILLER_185_310 ();
 sky130_fd_sc_hs__fill_8 FILLER_185_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_185_326 ();
 sky130_fd_sc_hs__fill_8 FILLER_185_334 ();
 sky130_fd_sc_hs__fill_4 FILLER_185_342 ();
 sky130_fd_sc_hs__fill_2 FILLER_185_346 ();
 sky130_fd_sc_hs__fill_8 FILLER_185_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_185_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_185_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_185_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_185_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_185_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_185_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_185_405 ();
 sky130_fd_sc_hs__fill_1 FILLER_185_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_185_440 ();
 sky130_fd_sc_hs__fill_4 FILLER_185_448 ();
 sky130_fd_sc_hs__fill_4 FILLER_185_458 ();
 sky130_fd_sc_hs__fill_2 FILLER_185_462 ();
 sky130_fd_sc_hs__fill_8 FILLER_185_488 ();
 sky130_fd_sc_hs__fill_2 FILLER_185_496 ();
 sky130_fd_sc_hs__fill_8 FILLER_185_506 ();
 sky130_fd_sc_hs__fill_8 FILLER_185_514 ();
 sky130_fd_sc_hs__fill_8 FILLER_185_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_185_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_185_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_186_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_186_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_186_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_186_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_186_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_186_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_186_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_186_46 ();
 sky130_fd_sc_hs__fill_2 FILLER_186_54 ();
 sky130_fd_sc_hs__fill_1 FILLER_186_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_186_74 ();
 sky130_fd_sc_hs__fill_4 FILLER_186_82 ();
 sky130_fd_sc_hs__fill_1 FILLER_186_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_186_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_186_96 ();
 sky130_fd_sc_hs__fill_4 FILLER_186_104 ();
 sky130_fd_sc_hs__fill_2 FILLER_186_108 ();
 sky130_fd_sc_hs__fill_8 FILLER_186_116 ();
 sky130_fd_sc_hs__fill_8 FILLER_186_124 ();
 sky130_fd_sc_hs__fill_4 FILLER_186_132 ();
 sky130_fd_sc_hs__fill_1 FILLER_186_144 ();
 sky130_fd_sc_hs__fill_4 FILLER_186_146 ();
 sky130_fd_sc_hs__fill_2 FILLER_186_150 ();
 sky130_fd_sc_hs__fill_1 FILLER_186_152 ();
 sky130_fd_sc_hs__fill_8 FILLER_186_172 ();
 sky130_fd_sc_hs__fill_8 FILLER_186_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_186_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_186_220 ();
 sky130_fd_sc_hs__fill_4 FILLER_186_228 ();
 sky130_fd_sc_hs__fill_1 FILLER_186_232 ();
 sky130_fd_sc_hs__fill_2 FILLER_186_236 ();
 sky130_fd_sc_hs__fill_1 FILLER_186_238 ();
 sky130_fd_sc_hs__fill_2 FILLER_186_272 ();
 sky130_fd_sc_hs__fill_1 FILLER_186_274 ();
 sky130_fd_sc_hs__fill_4 FILLER_186_281 ();
 sky130_fd_sc_hs__fill_2 FILLER_186_285 ();
 sky130_fd_sc_hs__fill_8 FILLER_186_310 ();
 sky130_fd_sc_hs__fill_1 FILLER_186_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_186_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_186_328 ();
 sky130_fd_sc_hs__fill_4 FILLER_186_336 ();
 sky130_fd_sc_hs__fill_2 FILLER_186_340 ();
 sky130_fd_sc_hs__fill_1 FILLER_186_342 ();
 sky130_fd_sc_hs__fill_8 FILLER_186_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_186_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_186_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_186_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_186_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_186_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_186_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_186_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_186_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_186_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_186_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_186_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_186_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_186_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_186_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_186_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_186_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_186_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_186_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_186_494 ();
 sky130_fd_sc_hs__fill_4 FILLER_186_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_186_514 ();
 sky130_fd_sc_hs__fill_8 FILLER_186_522 ();
 sky130_fd_sc_hs__fill_8 FILLER_186_530 ();
 sky130_fd_sc_hs__fill_2 FILLER_186_538 ();
 sky130_fd_sc_hs__fill_8 FILLER_187_0 ();
 sky130_fd_sc_hs__fill_4 FILLER_187_8 ();
 sky130_fd_sc_hs__fill_1 FILLER_187_12 ();
 sky130_fd_sc_hs__fill_8 FILLER_187_21 ();
 sky130_fd_sc_hs__fill_8 FILLER_187_29 ();
 sky130_fd_sc_hs__fill_1 FILLER_187_37 ();
 sky130_fd_sc_hs__fill_1 FILLER_187_59 ();
 sky130_fd_sc_hs__fill_1 FILLER_187_75 ();
 sky130_fd_sc_hs__fill_4 FILLER_187_89 ();
 sky130_fd_sc_hs__fill_8 FILLER_187_117 ();
 sky130_fd_sc_hs__fill_4 FILLER_187_125 ();
 sky130_fd_sc_hs__fill_1 FILLER_187_129 ();
 sky130_fd_sc_hs__fill_8 FILLER_187_142 ();
 sky130_fd_sc_hs__fill_8 FILLER_187_150 ();
 sky130_fd_sc_hs__fill_4 FILLER_187_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_187_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_187_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_187_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_187_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_187_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_187_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_187_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_187_231 ();
 sky130_fd_sc_hs__fill_4 FILLER_187_277 ();
 sky130_fd_sc_hs__fill_8 FILLER_187_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_187_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_187_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_187_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_187_323 ();
 sky130_fd_sc_hs__fill_4 FILLER_187_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_187_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_187_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_187_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_187_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_187_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_187_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_187_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_187_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_187_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_187_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_187_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_187_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_187_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_187_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_187_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_187_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_187_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_187_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_187_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_187_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_187_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_187_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_187_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_187_521 ();
 sky130_fd_sc_hs__fill_4 FILLER_187_523 ();
 sky130_fd_sc_hs__fill_1 FILLER_187_527 ();
 sky130_fd_sc_hs__fill_4 FILLER_187_536 ();
 sky130_fd_sc_hs__fill_4 FILLER_188_0 ();
 sky130_fd_sc_hs__fill_1 FILLER_188_4 ();
 sky130_fd_sc_hs__fill_8 FILLER_188_13 ();
 sky130_fd_sc_hs__fill_8 FILLER_188_21 ();
 sky130_fd_sc_hs__fill_8 FILLER_188_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_188_38 ();
 sky130_fd_sc_hs__fill_4 FILLER_188_53 ();
 sky130_fd_sc_hs__fill_1 FILLER_188_57 ();
 sky130_fd_sc_hs__fill_2 FILLER_188_68 ();
 sky130_fd_sc_hs__fill_8 FILLER_188_77 ();
 sky130_fd_sc_hs__fill_2 FILLER_188_85 ();
 sky130_fd_sc_hs__fill_8 FILLER_188_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_188_96 ();
 sky130_fd_sc_hs__fill_2 FILLER_188_104 ();
 sky130_fd_sc_hs__fill_1 FILLER_188_106 ();
 sky130_fd_sc_hs__fill_8 FILLER_188_114 ();
 sky130_fd_sc_hs__fill_4 FILLER_188_122 ();
 sky130_fd_sc_hs__fill_2 FILLER_188_126 ();
 sky130_fd_sc_hs__fill_1 FILLER_188_128 ();
 sky130_fd_sc_hs__fill_4 FILLER_188_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_188_156 ();
 sky130_fd_sc_hs__fill_4 FILLER_188_164 ();
 sky130_fd_sc_hs__fill_8 FILLER_188_174 ();
 sky130_fd_sc_hs__fill_8 FILLER_188_182 ();
 sky130_fd_sc_hs__fill_4 FILLER_188_190 ();
 sky130_fd_sc_hs__fill_2 FILLER_188_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_188_196 ();
 sky130_fd_sc_hs__fill_8 FILLER_188_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_188_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_188_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_188_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_188_236 ();
 sky130_fd_sc_hs__fill_2 FILLER_188_244 ();
 sky130_fd_sc_hs__fill_2 FILLER_188_249 ();
 sky130_fd_sc_hs__fill_2 FILLER_188_259 ();
 sky130_fd_sc_hs__fill_8 FILLER_188_262 ();
 sky130_fd_sc_hs__fill_4 FILLER_188_270 ();
 sky130_fd_sc_hs__fill_2 FILLER_188_274 ();
 sky130_fd_sc_hs__fill_8 FILLER_188_285 ();
 sky130_fd_sc_hs__fill_1 FILLER_188_293 ();
 sky130_fd_sc_hs__fill_8 FILLER_188_302 ();
 sky130_fd_sc_hs__fill_8 FILLER_188_310 ();
 sky130_fd_sc_hs__fill_1 FILLER_188_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_188_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_188_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_188_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_188_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_188_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_188_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_188_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_188_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_188_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_188_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_188_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_188_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_188_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_188_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_188_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_188_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_188_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_188_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_188_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_188_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_188_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_188_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_188_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_188_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_188_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_188_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_188_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_188_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_188_526 ();
 sky130_fd_sc_hs__fill_4 FILLER_188_534 ();
 sky130_fd_sc_hs__fill_2 FILLER_188_538 ();
 sky130_fd_sc_hs__fill_8 FILLER_189_0 ();
 sky130_fd_sc_hs__fill_4 FILLER_189_8 ();
 sky130_fd_sc_hs__fill_1 FILLER_189_12 ();
 sky130_fd_sc_hs__fill_8 FILLER_189_21 ();
 sky130_fd_sc_hs__fill_8 FILLER_189_29 ();
 sky130_fd_sc_hs__fill_8 FILLER_189_37 ();
 sky130_fd_sc_hs__fill_8 FILLER_189_45 ();
 sky130_fd_sc_hs__fill_2 FILLER_189_53 ();
 sky130_fd_sc_hs__fill_2 FILLER_189_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_189_71 ();
 sky130_fd_sc_hs__fill_8 FILLER_189_79 ();
 sky130_fd_sc_hs__fill_4 FILLER_189_87 ();
 sky130_fd_sc_hs__fill_1 FILLER_189_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_189_102 ();
 sky130_fd_sc_hs__fill_1 FILLER_189_110 ();
 sky130_fd_sc_hs__fill_8 FILLER_189_117 ();
 sky130_fd_sc_hs__fill_1 FILLER_189_125 ();
 sky130_fd_sc_hs__fill_1 FILLER_189_161 ();
 sky130_fd_sc_hs__fill_8 FILLER_189_166 ();
 sky130_fd_sc_hs__fill_8 FILLER_189_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_189_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_189_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_189_199 ();
 sky130_fd_sc_hs__fill_2 FILLER_189_207 ();
 sky130_fd_sc_hs__fill_1 FILLER_189_209 ();
 sky130_fd_sc_hs__fill_2 FILLER_189_215 ();
 sky130_fd_sc_hs__fill_1 FILLER_189_217 ();
 sky130_fd_sc_hs__fill_4 FILLER_189_227 ();
 sky130_fd_sc_hs__fill_1 FILLER_189_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_189_233 ();
 sky130_fd_sc_hs__fill_2 FILLER_189_241 ();
 sky130_fd_sc_hs__fill_2 FILLER_189_250 ();
 sky130_fd_sc_hs__fill_8 FILLER_189_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_189_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_189_291 ();
 sky130_fd_sc_hs__fill_2 FILLER_189_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_189_313 ();
 sky130_fd_sc_hs__fill_4 FILLER_189_321 ();
 sky130_fd_sc_hs__fill_2 FILLER_189_345 ();
 sky130_fd_sc_hs__fill_1 FILLER_189_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_189_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_189_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_189_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_189_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_189_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_189_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_189_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_189_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_189_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_189_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_189_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_189_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_189_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_189_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_189_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_189_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_189_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_189_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_189_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_189_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_189_497 ();
 sky130_fd_sc_hs__fill_1 FILLER_189_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_189_514 ();
 sky130_fd_sc_hs__fill_8 FILLER_189_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_189_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_189_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_190_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_190_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_190_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_190_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_190_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_190_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_190_38 ();
 sky130_fd_sc_hs__fill_4 FILLER_190_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_190_69 ();
 sky130_fd_sc_hs__fill_8 FILLER_190_77 ();
 sky130_fd_sc_hs__fill_2 FILLER_190_85 ();
 sky130_fd_sc_hs__fill_1 FILLER_190_88 ();
 sky130_fd_sc_hs__fill_4 FILLER_190_99 ();
 sky130_fd_sc_hs__fill_1 FILLER_190_103 ();
 sky130_fd_sc_hs__fill_8 FILLER_190_110 ();
 sky130_fd_sc_hs__fill_8 FILLER_190_118 ();
 sky130_fd_sc_hs__fill_8 FILLER_190_126 ();
 sky130_fd_sc_hs__fill_8 FILLER_190_134 ();
 sky130_fd_sc_hs__fill_2 FILLER_190_142 ();
 sky130_fd_sc_hs__fill_1 FILLER_190_144 ();
 sky130_fd_sc_hs__fill_4 FILLER_190_146 ();
 sky130_fd_sc_hs__fill_2 FILLER_190_150 ();
 sky130_fd_sc_hs__fill_1 FILLER_190_152 ();
 sky130_fd_sc_hs__fill_4 FILLER_190_171 ();
 sky130_fd_sc_hs__fill_4 FILLER_190_189 ();
 sky130_fd_sc_hs__fill_2 FILLER_190_193 ();
 sky130_fd_sc_hs__fill_4 FILLER_190_198 ();
 sky130_fd_sc_hs__fill_1 FILLER_190_202 ();
 sky130_fd_sc_hs__fill_4 FILLER_190_218 ();
 sky130_fd_sc_hs__fill_8 FILLER_190_229 ();
 sky130_fd_sc_hs__fill_2 FILLER_190_237 ();
 sky130_fd_sc_hs__fill_1 FILLER_190_239 ();
 sky130_fd_sc_hs__fill_8 FILLER_190_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_190_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_190_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_190_286 ();
 sky130_fd_sc_hs__fill_1 FILLER_190_294 ();
 sky130_fd_sc_hs__fill_4 FILLER_190_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_190_332 ();
 sky130_fd_sc_hs__fill_8 FILLER_190_340 ();
 sky130_fd_sc_hs__fill_8 FILLER_190_348 ();
 sky130_fd_sc_hs__fill_8 FILLER_190_356 ();
 sky130_fd_sc_hs__fill_8 FILLER_190_364 ();
 sky130_fd_sc_hs__fill_4 FILLER_190_372 ();
 sky130_fd_sc_hs__fill_1 FILLER_190_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_190_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_190_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_190_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_190_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_190_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_190_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_190_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_190_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_190_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_190_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_190_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_190_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_190_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_190_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_190_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_190_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_190_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_190_502 ();
 sky130_fd_sc_hs__fill_2 FILLER_190_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_190_520 ();
 sky130_fd_sc_hs__fill_8 FILLER_190_528 ();
 sky130_fd_sc_hs__fill_4 FILLER_190_536 ();
 sky130_fd_sc_hs__fill_8 FILLER_191_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_191_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_191_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_191_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_191_37 ();
 sky130_fd_sc_hs__fill_8 FILLER_191_45 ();
 sky130_fd_sc_hs__fill_4 FILLER_191_53 ();
 sky130_fd_sc_hs__fill_1 FILLER_191_57 ();
 sky130_fd_sc_hs__fill_8 FILLER_191_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_191_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_191_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_191_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_191_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_191_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_191_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_191_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_191_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_191_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_191_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_191_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_191_149 ();
 sky130_fd_sc_hs__fill_4 FILLER_191_160 ();
 sky130_fd_sc_hs__fill_4 FILLER_191_167 ();
 sky130_fd_sc_hs__fill_4 FILLER_191_185 ();
 sky130_fd_sc_hs__fill_1 FILLER_191_189 ();
 sky130_fd_sc_hs__fill_8 FILLER_191_200 ();
 sky130_fd_sc_hs__fill_1 FILLER_191_208 ();
 sky130_fd_sc_hs__fill_4 FILLER_191_226 ();
 sky130_fd_sc_hs__fill_2 FILLER_191_230 ();
 sky130_fd_sc_hs__fill_8 FILLER_191_233 ();
 sky130_fd_sc_hs__fill_2 FILLER_191_241 ();
 sky130_fd_sc_hs__fill_4 FILLER_191_267 ();
 sky130_fd_sc_hs__fill_2 FILLER_191_271 ();
 sky130_fd_sc_hs__fill_1 FILLER_191_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_191_278 ();
 sky130_fd_sc_hs__fill_1 FILLER_191_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_191_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_191_299 ();
 sky130_fd_sc_hs__fill_4 FILLER_191_307 ();
 sky130_fd_sc_hs__fill_2 FILLER_191_311 ();
 sky130_fd_sc_hs__fill_1 FILLER_191_313 ();
 sky130_fd_sc_hs__fill_8 FILLER_191_326 ();
 sky130_fd_sc_hs__fill_8 FILLER_191_334 ();
 sky130_fd_sc_hs__fill_4 FILLER_191_342 ();
 sky130_fd_sc_hs__fill_2 FILLER_191_346 ();
 sky130_fd_sc_hs__fill_8 FILLER_191_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_191_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_191_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_191_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_191_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_191_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_191_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_191_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_191_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_191_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_191_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_191_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_191_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_191_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_191_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_191_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_191_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_191_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_191_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_191_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_191_497 ();
 sky130_fd_sc_hs__fill_1 FILLER_191_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_191_514 ();
 sky130_fd_sc_hs__fill_8 FILLER_191_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_191_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_191_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_192_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_192_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_30 ();
 sky130_fd_sc_hs__fill_2 FILLER_192_38 ();
 sky130_fd_sc_hs__fill_1 FILLER_192_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_67 ();
 sky130_fd_sc_hs__fill_2 FILLER_192_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_192_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_178 ();
 sky130_fd_sc_hs__fill_4 FILLER_192_186 ();
 sky130_fd_sc_hs__fill_2 FILLER_192_190 ();
 sky130_fd_sc_hs__fill_1 FILLER_192_192 ();
 sky130_fd_sc_hs__fill_4 FILLER_192_196 ();
 sky130_fd_sc_hs__fill_2 FILLER_192_200 ();
 sky130_fd_sc_hs__fill_1 FILLER_192_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_204 ();
 sky130_fd_sc_hs__fill_2 FILLER_192_212 ();
 sky130_fd_sc_hs__fill_1 FILLER_192_214 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_192_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_262 ();
 sky130_fd_sc_hs__fill_4 FILLER_192_270 ();
 sky130_fd_sc_hs__fill_1 FILLER_192_274 ();
 sky130_fd_sc_hs__fill_1 FILLER_192_280 ();
 sky130_fd_sc_hs__fill_4 FILLER_192_289 ();
 sky130_fd_sc_hs__fill_1 FILLER_192_293 ();
 sky130_fd_sc_hs__fill_1 FILLER_192_302 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_308 ();
 sky130_fd_sc_hs__fill_2 FILLER_192_316 ();
 sky130_fd_sc_hs__fill_1 FILLER_192_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_192_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_192_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_192_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_192_526 ();
 sky130_fd_sc_hs__fill_4 FILLER_192_534 ();
 sky130_fd_sc_hs__fill_2 FILLER_192_538 ();
 sky130_fd_sc_hs__fill_8 FILLER_193_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_193_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_193_16 ();
 sky130_fd_sc_hs__fill_1 FILLER_193_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_193_33 ();
 sky130_fd_sc_hs__fill_2 FILLER_193_53 ();
 sky130_fd_sc_hs__fill_8 FILLER_193_59 ();
 sky130_fd_sc_hs__fill_2 FILLER_193_70 ();
 sky130_fd_sc_hs__fill_1 FILLER_193_72 ();
 sky130_fd_sc_hs__fill_8 FILLER_193_78 ();
 sky130_fd_sc_hs__fill_2 FILLER_193_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_193_100 ();
 sky130_fd_sc_hs__fill_8 FILLER_193_108 ();
 sky130_fd_sc_hs__fill_8 FILLER_193_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_193_125 ();
 sky130_fd_sc_hs__fill_1 FILLER_193_133 ();
 sky130_fd_sc_hs__fill_4 FILLER_193_169 ();
 sky130_fd_sc_hs__fill_1 FILLER_193_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_193_175 ();
 sky130_fd_sc_hs__fill_1 FILLER_193_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_193_205 ();
 sky130_fd_sc_hs__fill_8 FILLER_193_213 ();
 sky130_fd_sc_hs__fill_8 FILLER_193_221 ();
 sky130_fd_sc_hs__fill_2 FILLER_193_229 ();
 sky130_fd_sc_hs__fill_1 FILLER_193_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_193_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_193_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_193_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_193_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_193_265 ();
 sky130_fd_sc_hs__fill_4 FILLER_193_273 ();
 sky130_fd_sc_hs__fill_1 FILLER_193_277 ();
 sky130_fd_sc_hs__fill_4 FILLER_193_291 ();
 sky130_fd_sc_hs__fill_1 FILLER_193_295 ();
 sky130_fd_sc_hs__fill_1 FILLER_193_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_193_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_193_336 ();
 sky130_fd_sc_hs__fill_4 FILLER_193_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_193_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_193_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_193_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_193_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_193_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_193_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_193_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_193_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_193_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_193_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_193_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_193_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_193_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_193_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_193_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_193_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_193_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_193_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_193_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_193_489 ();
 sky130_fd_sc_hs__fill_1 FILLER_193_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_193_506 ();
 sky130_fd_sc_hs__fill_8 FILLER_193_514 ();
 sky130_fd_sc_hs__fill_8 FILLER_193_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_193_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_193_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_194_0 ();
 sky130_fd_sc_hs__fill_4 FILLER_194_8 ();
 sky130_fd_sc_hs__fill_1 FILLER_194_12 ();
 sky130_fd_sc_hs__fill_8 FILLER_194_21 ();
 sky130_fd_sc_hs__fill_4 FILLER_194_30 ();
 sky130_fd_sc_hs__fill_1 FILLER_194_34 ();
 sky130_fd_sc_hs__fill_8 FILLER_194_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_194_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_194_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_194_108 ();
 sky130_fd_sc_hs__fill_8 FILLER_194_116 ();
 sky130_fd_sc_hs__fill_8 FILLER_194_124 ();
 sky130_fd_sc_hs__fill_1 FILLER_194_132 ();
 sky130_fd_sc_hs__fill_8 FILLER_194_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_194_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_194_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_194_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_194_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_194_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_194_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_194_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_194_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_194_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_194_220 ();
 sky130_fd_sc_hs__fill_4 FILLER_194_228 ();
 sky130_fd_sc_hs__fill_4 FILLER_194_244 ();
 sky130_fd_sc_hs__fill_1 FILLER_194_248 ();
 sky130_fd_sc_hs__fill_4 FILLER_194_262 ();
 sky130_fd_sc_hs__fill_2 FILLER_194_266 ();
 sky130_fd_sc_hs__fill_1 FILLER_194_280 ();
 sky130_fd_sc_hs__fill_8 FILLER_194_292 ();
 sky130_fd_sc_hs__fill_8 FILLER_194_300 ();
 sky130_fd_sc_hs__fill_8 FILLER_194_308 ();
 sky130_fd_sc_hs__fill_2 FILLER_194_316 ();
 sky130_fd_sc_hs__fill_1 FILLER_194_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_194_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_194_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_194_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_194_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_194_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_194_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_194_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_194_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_194_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_194_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_194_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_194_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_194_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_194_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_194_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_194_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_194_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_194_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_194_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_194_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_194_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_194_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_194_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_194_492 ();
 sky130_fd_sc_hs__fill_4 FILLER_194_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_194_506 ();
 sky130_fd_sc_hs__fill_8 FILLER_194_514 ();
 sky130_fd_sc_hs__fill_8 FILLER_194_522 ();
 sky130_fd_sc_hs__fill_8 FILLER_194_530 ();
 sky130_fd_sc_hs__fill_2 FILLER_194_538 ();
 sky130_fd_sc_hs__fill_4 FILLER_195_0 ();
 sky130_fd_sc_hs__fill_1 FILLER_195_4 ();
 sky130_fd_sc_hs__fill_1 FILLER_195_13 ();
 sky130_fd_sc_hs__fill_2 FILLER_195_23 ();
 sky130_fd_sc_hs__fill_1 FILLER_195_25 ();
 sky130_fd_sc_hs__fill_1 FILLER_195_57 ();
 sky130_fd_sc_hs__fill_2 FILLER_195_59 ();
 sky130_fd_sc_hs__fill_1 FILLER_195_61 ();
 sky130_fd_sc_hs__fill_8 FILLER_195_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_195_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_195_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_195_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_195_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_195_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_195_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_195_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_195_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_195_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_195_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_195_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_195_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_195_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_195_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_195_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_195_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_195_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_195_249 ();
 sky130_fd_sc_hs__fill_4 FILLER_195_257 ();
 sky130_fd_sc_hs__fill_2 FILLER_195_261 ();
 sky130_fd_sc_hs__fill_4 FILLER_195_284 ();
 sky130_fd_sc_hs__fill_2 FILLER_195_288 ();
 sky130_fd_sc_hs__fill_8 FILLER_195_302 ();
 sky130_fd_sc_hs__fill_8 FILLER_195_310 ();
 sky130_fd_sc_hs__fill_8 FILLER_195_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_195_326 ();
 sky130_fd_sc_hs__fill_8 FILLER_195_334 ();
 sky130_fd_sc_hs__fill_4 FILLER_195_342 ();
 sky130_fd_sc_hs__fill_2 FILLER_195_346 ();
 sky130_fd_sc_hs__fill_8 FILLER_195_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_195_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_195_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_195_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_195_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_195_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_195_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_195_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_195_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_195_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_195_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_195_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_195_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_195_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_195_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_195_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_195_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_195_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_195_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_195_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_195_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_195_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_195_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_195_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_195_523 ();
 sky130_fd_sc_hs__fill_1 FILLER_195_531 ();
 sky130_fd_sc_hs__fill_8 FILLER_196_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_196_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_196_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_196_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_196_28 ();
 sky130_fd_sc_hs__fill_1 FILLER_196_30 ();
 sky130_fd_sc_hs__fill_4 FILLER_196_38 ();
 sky130_fd_sc_hs__fill_2 FILLER_196_42 ();
 sky130_fd_sc_hs__fill_4 FILLER_196_82 ();
 sky130_fd_sc_hs__fill_1 FILLER_196_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_196_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_196_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_196_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_196_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_196_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_196_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_196_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_196_144 ();
 sky130_fd_sc_hs__fill_2 FILLER_196_146 ();
 sky130_fd_sc_hs__fill_1 FILLER_196_148 ();
 sky130_fd_sc_hs__fill_8 FILLER_196_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_196_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_196_239 ();
 sky130_fd_sc_hs__fill_8 FILLER_196_247 ();
 sky130_fd_sc_hs__fill_4 FILLER_196_255 ();
 sky130_fd_sc_hs__fill_2 FILLER_196_259 ();
 sky130_fd_sc_hs__fill_8 FILLER_196_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_196_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_196_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_196_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_196_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_196_302 ();
 sky130_fd_sc_hs__fill_8 FILLER_196_310 ();
 sky130_fd_sc_hs__fill_1 FILLER_196_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_196_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_196_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_196_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_196_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_196_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_196_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_196_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_196_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_196_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_196_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_196_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_196_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_196_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_196_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_196_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_196_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_196_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_196_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_196_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_196_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_196_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_196_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_196_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_196_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_196_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_196_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_196_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_196_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_196_526 ();
 sky130_fd_sc_hs__fill_4 FILLER_196_534 ();
 sky130_fd_sc_hs__fill_2 FILLER_196_538 ();
 sky130_fd_sc_hs__fill_4 FILLER_197_0 ();
 sky130_fd_sc_hs__fill_1 FILLER_197_4 ();
 sky130_fd_sc_hs__fill_8 FILLER_197_13 ();
 sky130_fd_sc_hs__fill_8 FILLER_197_21 ();
 sky130_fd_sc_hs__fill_8 FILLER_197_29 ();
 sky130_fd_sc_hs__fill_8 FILLER_197_37 ();
 sky130_fd_sc_hs__fill_8 FILLER_197_45 ();
 sky130_fd_sc_hs__fill_4 FILLER_197_53 ();
 sky130_fd_sc_hs__fill_1 FILLER_197_57 ();
 sky130_fd_sc_hs__fill_2 FILLER_197_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_197_80 ();
 sky130_fd_sc_hs__fill_8 FILLER_197_117 ();
 sky130_fd_sc_hs__fill_4 FILLER_197_125 ();
 sky130_fd_sc_hs__fill_2 FILLER_197_129 ();
 sky130_fd_sc_hs__fill_1 FILLER_197_131 ();
 sky130_fd_sc_hs__fill_4 FILLER_197_167 ();
 sky130_fd_sc_hs__fill_2 FILLER_197_171 ();
 sky130_fd_sc_hs__fill_1 FILLER_197_173 ();
 sky130_fd_sc_hs__fill_4 FILLER_197_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_197_214 ();
 sky130_fd_sc_hs__fill_2 FILLER_197_222 ();
 sky130_fd_sc_hs__fill_1 FILLER_197_224 ();
 sky130_fd_sc_hs__fill_4 FILLER_197_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_197_233 ();
 sky130_fd_sc_hs__fill_4 FILLER_197_241 ();
 sky130_fd_sc_hs__fill_2 FILLER_197_258 ();
 sky130_fd_sc_hs__fill_1 FILLER_197_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_197_274 ();
 sky130_fd_sc_hs__fill_8 FILLER_197_282 ();
 sky130_fd_sc_hs__fill_4 FILLER_197_291 ();
 sky130_fd_sc_hs__fill_2 FILLER_197_295 ();
 sky130_fd_sc_hs__fill_8 FILLER_197_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_197_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_197_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_197_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_197_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_197_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_197_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_197_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_197_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_197_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_197_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_197_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_197_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_197_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_197_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_197_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_197_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_197_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_197_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_197_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_197_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_197_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_197_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_197_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_197_489 ();
 sky130_fd_sc_hs__fill_1 FILLER_197_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_197_506 ();
 sky130_fd_sc_hs__fill_8 FILLER_197_514 ();
 sky130_fd_sc_hs__fill_8 FILLER_197_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_197_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_197_539 ();
 sky130_fd_sc_hs__fill_2 FILLER_198_0 ();
 sky130_fd_sc_hs__fill_1 FILLER_198_2 ();
 sky130_fd_sc_hs__fill_8 FILLER_198_11 ();
 sky130_fd_sc_hs__fill_8 FILLER_198_19 ();
 sky130_fd_sc_hs__fill_2 FILLER_198_27 ();
 sky130_fd_sc_hs__fill_8 FILLER_198_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_198_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_198_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_198_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_198_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_198_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_198_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_198_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_198_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_198_96 ();
 sky130_fd_sc_hs__fill_4 FILLER_198_104 ();
 sky130_fd_sc_hs__fill_2 FILLER_198_108 ();
 sky130_fd_sc_hs__fill_8 FILLER_198_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_198_154 ();
 sky130_fd_sc_hs__fill_4 FILLER_198_162 ();
 sky130_fd_sc_hs__fill_2 FILLER_198_166 ();
 sky130_fd_sc_hs__fill_4 FILLER_198_204 ();
 sky130_fd_sc_hs__fill_1 FILLER_198_220 ();
 sky130_fd_sc_hs__fill_4 FILLER_198_240 ();
 sky130_fd_sc_hs__fill_4 FILLER_198_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_198_275 ();
 sky130_fd_sc_hs__fill_8 FILLER_198_283 ();
 sky130_fd_sc_hs__fill_4 FILLER_198_291 ();
 sky130_fd_sc_hs__fill_2 FILLER_198_295 ();
 sky130_fd_sc_hs__fill_4 FILLER_198_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_198_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_198_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_198_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_198_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_198_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_198_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_198_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_198_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_198_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_198_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_198_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_198_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_198_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_198_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_198_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_198_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_198_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_198_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_198_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_198_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_198_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_198_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_198_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_198_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_198_494 ();
 sky130_fd_sc_hs__fill_4 FILLER_198_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_198_514 ();
 sky130_fd_sc_hs__fill_8 FILLER_198_522 ();
 sky130_fd_sc_hs__fill_8 FILLER_198_530 ();
 sky130_fd_sc_hs__fill_2 FILLER_198_538 ();
 sky130_fd_sc_hs__fill_8 FILLER_199_0 ();
 sky130_fd_sc_hs__fill_4 FILLER_199_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_199_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_199_32 ();
 sky130_fd_sc_hs__fill_8 FILLER_199_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_199_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_199_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_199_59 ();
 sky130_fd_sc_hs__fill_1 FILLER_199_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_199_71 ();
 sky130_fd_sc_hs__fill_8 FILLER_199_79 ();
 sky130_fd_sc_hs__fill_4 FILLER_199_87 ();
 sky130_fd_sc_hs__fill_2 FILLER_199_91 ();
 sky130_fd_sc_hs__fill_1 FILLER_199_93 ();
 sky130_fd_sc_hs__fill_1 FILLER_199_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_199_153 ();
 sky130_fd_sc_hs__fill_8 FILLER_199_161 ();
 sky130_fd_sc_hs__fill_4 FILLER_199_169 ();
 sky130_fd_sc_hs__fill_1 FILLER_199_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_199_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_199_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_199_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_199_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_199_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_199_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_199_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_199_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_199_233 ();
 sky130_fd_sc_hs__fill_4 FILLER_199_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_199_279 ();
 sky130_fd_sc_hs__fill_2 FILLER_199_287 ();
 sky130_fd_sc_hs__fill_1 FILLER_199_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_199_291 ();
 sky130_fd_sc_hs__fill_1 FILLER_199_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_199_313 ();
 sky130_fd_sc_hs__fill_8 FILLER_199_321 ();
 sky130_fd_sc_hs__fill_8 FILLER_199_329 ();
 sky130_fd_sc_hs__fill_8 FILLER_199_337 ();
 sky130_fd_sc_hs__fill_2 FILLER_199_345 ();
 sky130_fd_sc_hs__fill_1 FILLER_199_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_199_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_199_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_199_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_199_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_199_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_199_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_199_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_199_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_199_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_199_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_199_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_199_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_199_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_199_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_199_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_199_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_199_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_199_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_199_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_199_489 ();
 sky130_fd_sc_hs__fill_1 FILLER_199_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_199_506 ();
 sky130_fd_sc_hs__fill_8 FILLER_199_514 ();
 sky130_fd_sc_hs__fill_8 FILLER_199_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_199_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_199_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_200_0 ();
 sky130_fd_sc_hs__fill_4 FILLER_200_8 ();
 sky130_fd_sc_hs__fill_2 FILLER_200_12 ();
 sky130_fd_sc_hs__fill_8 FILLER_200_39 ();
 sky130_fd_sc_hs__fill_8 FILLER_200_47 ();
 sky130_fd_sc_hs__fill_8 FILLER_200_55 ();
 sky130_fd_sc_hs__fill_8 FILLER_200_63 ();
 sky130_fd_sc_hs__fill_8 FILLER_200_71 ();
 sky130_fd_sc_hs__fill_8 FILLER_200_79 ();
 sky130_fd_sc_hs__fill_2 FILLER_200_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_200_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_200_133 ();
 sky130_fd_sc_hs__fill_4 FILLER_200_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_200_146 ();
 sky130_fd_sc_hs__fill_2 FILLER_200_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_200_191 ();
 sky130_fd_sc_hs__fill_4 FILLER_200_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_200_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_200_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_200_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_200_228 ();
 sky130_fd_sc_hs__fill_4 FILLER_200_236 ();
 sky130_fd_sc_hs__fill_4 FILLER_200_262 ();
 sky130_fd_sc_hs__fill_1 FILLER_200_266 ();
 sky130_fd_sc_hs__fill_8 FILLER_200_279 ();
 sky130_fd_sc_hs__fill_4 FILLER_200_287 ();
 sky130_fd_sc_hs__fill_2 FILLER_200_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_200_306 ();
 sky130_fd_sc_hs__fill_4 FILLER_200_314 ();
 sky130_fd_sc_hs__fill_1 FILLER_200_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_200_340 ();
 sky130_fd_sc_hs__fill_8 FILLER_200_348 ();
 sky130_fd_sc_hs__fill_8 FILLER_200_356 ();
 sky130_fd_sc_hs__fill_8 FILLER_200_364 ();
 sky130_fd_sc_hs__fill_4 FILLER_200_372 ();
 sky130_fd_sc_hs__fill_1 FILLER_200_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_200_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_200_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_200_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_200_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_200_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_200_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_200_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_200_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_200_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_200_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_200_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_200_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_200_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_200_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_200_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_200_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_200_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_200_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_200_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_200_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_200_526 ();
 sky130_fd_sc_hs__fill_4 FILLER_200_534 ();
 sky130_fd_sc_hs__fill_2 FILLER_200_538 ();
 sky130_fd_sc_hs__fill_8 FILLER_201_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_201_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_201_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_201_24 ();
 sky130_fd_sc_hs__fill_8 FILLER_201_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_201_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_201_59 ();
 sky130_fd_sc_hs__fill_2 FILLER_201_71 ();
 sky130_fd_sc_hs__fill_1 FILLER_201_73 ();
 sky130_fd_sc_hs__fill_8 FILLER_201_82 ();
 sky130_fd_sc_hs__fill_8 FILLER_201_90 ();
 sky130_fd_sc_hs__fill_8 FILLER_201_98 ();
 sky130_fd_sc_hs__fill_8 FILLER_201_106 ();
 sky130_fd_sc_hs__fill_2 FILLER_201_114 ();
 sky130_fd_sc_hs__fill_1 FILLER_201_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_201_153 ();
 sky130_fd_sc_hs__fill_8 FILLER_201_161 ();
 sky130_fd_sc_hs__fill_4 FILLER_201_169 ();
 sky130_fd_sc_hs__fill_1 FILLER_201_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_201_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_201_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_201_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_201_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_201_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_201_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_201_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_201_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_201_233 ();
 sky130_fd_sc_hs__fill_4 FILLER_201_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_201_258 ();
 sky130_fd_sc_hs__fill_8 FILLER_201_266 ();
 sky130_fd_sc_hs__fill_8 FILLER_201_274 ();
 sky130_fd_sc_hs__fill_2 FILLER_201_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_201_305 ();
 sky130_fd_sc_hs__fill_8 FILLER_201_313 ();
 sky130_fd_sc_hs__fill_8 FILLER_201_321 ();
 sky130_fd_sc_hs__fill_8 FILLER_201_329 ();
 sky130_fd_sc_hs__fill_8 FILLER_201_337 ();
 sky130_fd_sc_hs__fill_2 FILLER_201_345 ();
 sky130_fd_sc_hs__fill_1 FILLER_201_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_201_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_201_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_201_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_201_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_201_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_201_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_201_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_201_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_201_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_201_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_201_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_201_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_201_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_201_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_201_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_201_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_201_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_201_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_201_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_201_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_201_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_201_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_201_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_201_521 ();
 sky130_fd_sc_hs__fill_4 FILLER_201_523 ();
 sky130_fd_sc_hs__fill_1 FILLER_201_527 ();
 sky130_fd_sc_hs__fill_4 FILLER_201_536 ();
 sky130_fd_sc_hs__fill_4 FILLER_202_0 ();
 sky130_fd_sc_hs__fill_1 FILLER_202_4 ();
 sky130_fd_sc_hs__fill_8 FILLER_202_30 ();
 sky130_fd_sc_hs__fill_2 FILLER_202_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_202_77 ();
 sky130_fd_sc_hs__fill_2 FILLER_202_85 ();
 sky130_fd_sc_hs__fill_8 FILLER_202_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_202_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_202_107 ();
 sky130_fd_sc_hs__fill_8 FILLER_202_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_202_123 ();
 sky130_fd_sc_hs__fill_8 FILLER_202_131 ();
 sky130_fd_sc_hs__fill_4 FILLER_202_139 ();
 sky130_fd_sc_hs__fill_2 FILLER_202_143 ();
 sky130_fd_sc_hs__fill_8 FILLER_202_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_202_154 ();
 sky130_fd_sc_hs__fill_2 FILLER_202_162 ();
 sky130_fd_sc_hs__fill_4 FILLER_202_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_202_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_202_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_202_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_202_228 ();
 sky130_fd_sc_hs__fill_4 FILLER_202_236 ();
 sky130_fd_sc_hs__fill_1 FILLER_202_240 ();
 sky130_fd_sc_hs__fill_4 FILLER_202_254 ();
 sky130_fd_sc_hs__fill_2 FILLER_202_258 ();
 sky130_fd_sc_hs__fill_1 FILLER_202_260 ();
 sky130_fd_sc_hs__fill_1 FILLER_202_262 ();
 sky130_fd_sc_hs__fill_4 FILLER_202_279 ();
 sky130_fd_sc_hs__fill_8 FILLER_202_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_202_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_202_307 ();
 sky130_fd_sc_hs__fill_4 FILLER_202_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_202_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_202_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_202_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_202_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_202_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_202_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_202_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_202_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_202_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_202_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_202_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_202_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_202_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_202_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_202_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_202_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_202_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_202_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_202_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_202_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_202_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_202_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_202_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_202_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_202_494 ();
 sky130_fd_sc_hs__fill_2 FILLER_202_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_202_512 ();
 sky130_fd_sc_hs__fill_8 FILLER_202_520 ();
 sky130_fd_sc_hs__fill_8 FILLER_202_528 ();
 sky130_fd_sc_hs__fill_4 FILLER_202_536 ();
 sky130_fd_sc_hs__fill_4 FILLER_203_0 ();
 sky130_fd_sc_hs__fill_2 FILLER_203_4 ();
 sky130_fd_sc_hs__fill_8 FILLER_203_14 ();
 sky130_fd_sc_hs__fill_2 FILLER_203_22 ();
 sky130_fd_sc_hs__fill_1 FILLER_203_24 ();
 sky130_fd_sc_hs__fill_4 FILLER_203_59 ();
 sky130_fd_sc_hs__fill_2 FILLER_203_63 ();
 sky130_fd_sc_hs__fill_1 FILLER_203_65 ();
 sky130_fd_sc_hs__fill_8 FILLER_203_101 ();
 sky130_fd_sc_hs__fill_4 FILLER_203_109 ();
 sky130_fd_sc_hs__fill_2 FILLER_203_113 ();
 sky130_fd_sc_hs__fill_1 FILLER_203_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_203_117 ();
 sky130_fd_sc_hs__fill_2 FILLER_203_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_203_162 ();
 sky130_fd_sc_hs__fill_4 FILLER_203_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_203_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_203_183 ();
 sky130_fd_sc_hs__fill_4 FILLER_203_191 ();
 sky130_fd_sc_hs__fill_2 FILLER_203_195 ();
 sky130_fd_sc_hs__fill_4 FILLER_203_218 ();
 sky130_fd_sc_hs__fill_2 FILLER_203_222 ();
 sky130_fd_sc_hs__fill_1 FILLER_203_231 ();
 sky130_fd_sc_hs__fill_4 FILLER_203_233 ();
 sky130_fd_sc_hs__fill_1 FILLER_203_237 ();
 sky130_fd_sc_hs__fill_8 FILLER_203_251 ();
 sky130_fd_sc_hs__fill_8 FILLER_203_259 ();
 sky130_fd_sc_hs__fill_8 FILLER_203_267 ();
 sky130_fd_sc_hs__fill_4 FILLER_203_275 ();
 sky130_fd_sc_hs__fill_2 FILLER_203_288 ();
 sky130_fd_sc_hs__fill_8 FILLER_203_325 ();
 sky130_fd_sc_hs__fill_8 FILLER_203_333 ();
 sky130_fd_sc_hs__fill_4 FILLER_203_341 ();
 sky130_fd_sc_hs__fill_2 FILLER_203_345 ();
 sky130_fd_sc_hs__fill_1 FILLER_203_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_203_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_203_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_203_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_203_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_203_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_203_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_203_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_203_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_203_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_203_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_203_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_203_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_203_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_203_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_203_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_203_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_203_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_203_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_203_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_203_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_203_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_203_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_203_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_203_521 ();
 sky130_fd_sc_hs__fill_2 FILLER_203_523 ();
 sky130_fd_sc_hs__fill_1 FILLER_203_525 ();
 sky130_fd_sc_hs__fill_4 FILLER_203_534 ();
 sky130_fd_sc_hs__fill_2 FILLER_203_538 ();
 sky130_fd_sc_hs__fill_8 FILLER_204_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_204_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_204_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_204_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_204_28 ();
 sky130_fd_sc_hs__fill_4 FILLER_204_30 ();
 sky130_fd_sc_hs__fill_1 FILLER_204_34 ();
 sky130_fd_sc_hs__fill_8 FILLER_204_52 ();
 sky130_fd_sc_hs__fill_4 FILLER_204_60 ();
 sky130_fd_sc_hs__fill_1 FILLER_204_64 ();
 sky130_fd_sc_hs__fill_4 FILLER_204_80 ();
 sky130_fd_sc_hs__fill_2 FILLER_204_84 ();
 sky130_fd_sc_hs__fill_1 FILLER_204_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_204_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_204_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_204_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_204_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_204_120 ();
 sky130_fd_sc_hs__fill_4 FILLER_204_128 ();
 sky130_fd_sc_hs__fill_1 FILLER_204_132 ();
 sky130_fd_sc_hs__fill_8 FILLER_204_146 ();
 sky130_fd_sc_hs__fill_4 FILLER_204_154 ();
 sky130_fd_sc_hs__fill_2 FILLER_204_158 ();
 sky130_fd_sc_hs__fill_8 FILLER_204_195 ();
 sky130_fd_sc_hs__fill_8 FILLER_204_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_204_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_204_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_204_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_204_236 ();
 sky130_fd_sc_hs__fill_8 FILLER_204_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_204_252 ();
 sky130_fd_sc_hs__fill_1 FILLER_204_260 ();
 sky130_fd_sc_hs__fill_2 FILLER_204_262 ();
 sky130_fd_sc_hs__fill_1 FILLER_204_264 ();
 sky130_fd_sc_hs__fill_8 FILLER_204_301 ();
 sky130_fd_sc_hs__fill_8 FILLER_204_309 ();
 sky130_fd_sc_hs__fill_2 FILLER_204_317 ();
 sky130_fd_sc_hs__fill_8 FILLER_204_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_204_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_204_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_204_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_204_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_204_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_204_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_204_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_204_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_204_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_204_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_204_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_204_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_204_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_204_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_204_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_204_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_204_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_204_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_204_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_204_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_204_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_204_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_204_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_204_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_204_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_204_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_204_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_204_526 ();
 sky130_fd_sc_hs__fill_4 FILLER_204_534 ();
 sky130_fd_sc_hs__fill_2 FILLER_204_538 ();
 sky130_fd_sc_hs__fill_8 FILLER_205_0 ();
 sky130_fd_sc_hs__fill_4 FILLER_205_8 ();
 sky130_fd_sc_hs__fill_1 FILLER_205_12 ();
 sky130_fd_sc_hs__fill_2 FILLER_205_21 ();
 sky130_fd_sc_hs__fill_1 FILLER_205_23 ();
 sky130_fd_sc_hs__fill_8 FILLER_205_46 ();
 sky130_fd_sc_hs__fill_4 FILLER_205_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_205_59 ();
 sky130_fd_sc_hs__fill_2 FILLER_205_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_205_82 ();
 sky130_fd_sc_hs__fill_8 FILLER_205_90 ();
 sky130_fd_sc_hs__fill_8 FILLER_205_98 ();
 sky130_fd_sc_hs__fill_8 FILLER_205_106 ();
 sky130_fd_sc_hs__fill_2 FILLER_205_114 ();
 sky130_fd_sc_hs__fill_4 FILLER_205_117 ();
 sky130_fd_sc_hs__fill_2 FILLER_205_121 ();
 sky130_fd_sc_hs__fill_8 FILLER_205_158 ();
 sky130_fd_sc_hs__fill_8 FILLER_205_166 ();
 sky130_fd_sc_hs__fill_8 FILLER_205_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_205_183 ();
 sky130_fd_sc_hs__fill_2 FILLER_205_191 ();
 sky130_fd_sc_hs__fill_1 FILLER_205_193 ();
 sky130_fd_sc_hs__fill_8 FILLER_205_215 ();
 sky130_fd_sc_hs__fill_8 FILLER_205_223 ();
 sky130_fd_sc_hs__fill_1 FILLER_205_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_205_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_205_241 ();
 sky130_fd_sc_hs__fill_1 FILLER_205_261 ();
 sky130_fd_sc_hs__fill_8 FILLER_205_267 ();
 sky130_fd_sc_hs__fill_8 FILLER_205_275 ();
 sky130_fd_sc_hs__fill_4 FILLER_205_283 ();
 sky130_fd_sc_hs__fill_2 FILLER_205_287 ();
 sky130_fd_sc_hs__fill_1 FILLER_205_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_205_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_205_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_205_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_205_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_205_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_205_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_205_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_205_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_205_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_205_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_205_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_205_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_205_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_205_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_205_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_205_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_205_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_205_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_205_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_205_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_205_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_205_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_205_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_205_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_205_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_205_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_205_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_205_489 ();
 sky130_fd_sc_hs__fill_1 FILLER_205_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_205_506 ();
 sky130_fd_sc_hs__fill_8 FILLER_205_514 ();
 sky130_fd_sc_hs__fill_8 FILLER_205_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_205_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_205_539 ();
 sky130_fd_sc_hs__fill_4 FILLER_206_0 ();
 sky130_fd_sc_hs__fill_2 FILLER_206_4 ();
 sky130_fd_sc_hs__fill_1 FILLER_206_6 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_15 ();
 sky130_fd_sc_hs__fill_4 FILLER_206_23 ();
 sky130_fd_sc_hs__fill_2 FILLER_206_27 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_43 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_51 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_75 ();
 sky130_fd_sc_hs__fill_4 FILLER_206_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_94 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_102 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_206_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_220 ();
 sky130_fd_sc_hs__fill_2 FILLER_206_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_253 ();
 sky130_fd_sc_hs__fill_2 FILLER_206_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_277 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_285 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_293 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_301 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_309 ();
 sky130_fd_sc_hs__fill_2 FILLER_206_317 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_206_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_206_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_206_492 ();
 sky130_fd_sc_hs__fill_4 FILLER_206_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_506 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_514 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_522 ();
 sky130_fd_sc_hs__fill_8 FILLER_206_530 ();
 sky130_fd_sc_hs__fill_2 FILLER_206_538 ();
 sky130_fd_sc_hs__fill_2 FILLER_207_0 ();
 sky130_fd_sc_hs__fill_2 FILLER_207_10 ();
 sky130_fd_sc_hs__fill_1 FILLER_207_12 ();
 sky130_fd_sc_hs__fill_4 FILLER_207_22 ();
 sky130_fd_sc_hs__fill_2 FILLER_207_26 ();
 sky130_fd_sc_hs__fill_1 FILLER_207_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_207_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_207_48 ();
 sky130_fd_sc_hs__fill_2 FILLER_207_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_207_59 ();
 sky130_fd_sc_hs__fill_1 FILLER_207_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_207_93 ();
 sky130_fd_sc_hs__fill_8 FILLER_207_101 ();
 sky130_fd_sc_hs__fill_4 FILLER_207_109 ();
 sky130_fd_sc_hs__fill_2 FILLER_207_113 ();
 sky130_fd_sc_hs__fill_1 FILLER_207_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_207_117 ();
 sky130_fd_sc_hs__fill_4 FILLER_207_125 ();
 sky130_fd_sc_hs__fill_1 FILLER_207_129 ();
 sky130_fd_sc_hs__fill_8 FILLER_207_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_207_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_207_175 ();
 sky130_fd_sc_hs__fill_2 FILLER_207_183 ();
 sky130_fd_sc_hs__fill_4 FILLER_207_206 ();
 sky130_fd_sc_hs__fill_1 FILLER_207_210 ();
 sky130_fd_sc_hs__fill_8 FILLER_207_254 ();
 sky130_fd_sc_hs__fill_8 FILLER_207_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_207_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_207_278 ();
 sky130_fd_sc_hs__fill_4 FILLER_207_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_207_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_207_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_207_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_207_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_207_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_207_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_207_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_207_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_207_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_207_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_207_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_207_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_207_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_207_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_207_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_207_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_207_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_207_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_207_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_207_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_207_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_207_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_207_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_207_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_207_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_207_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_207_481 ();
 sky130_fd_sc_hs__fill_4 FILLER_207_489 ();
 sky130_fd_sc_hs__fill_2 FILLER_207_493 ();
 sky130_fd_sc_hs__fill_1 FILLER_207_495 ();
 sky130_fd_sc_hs__fill_8 FILLER_207_506 ();
 sky130_fd_sc_hs__fill_8 FILLER_207_514 ();
 sky130_fd_sc_hs__fill_8 FILLER_207_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_207_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_207_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_208_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_208_8 ();
 sky130_fd_sc_hs__fill_1 FILLER_208_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_208_22 ();
 sky130_fd_sc_hs__fill_2 FILLER_208_26 ();
 sky130_fd_sc_hs__fill_1 FILLER_208_28 ();
 sky130_fd_sc_hs__fill_1 FILLER_208_33 ();
 sky130_fd_sc_hs__fill_4 FILLER_208_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_208_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_208_62 ();
 sky130_fd_sc_hs__fill_2 FILLER_208_70 ();
 sky130_fd_sc_hs__fill_1 FILLER_208_72 ();
 sky130_fd_sc_hs__fill_8 FILLER_208_77 ();
 sky130_fd_sc_hs__fill_2 FILLER_208_85 ();
 sky130_fd_sc_hs__fill_1 FILLER_208_94 ();
 sky130_fd_sc_hs__fill_1 FILLER_208_103 ();
 sky130_fd_sc_hs__fill_8 FILLER_208_122 ();
 sky130_fd_sc_hs__fill_2 FILLER_208_130 ();
 sky130_fd_sc_hs__fill_1 FILLER_208_132 ();
 sky130_fd_sc_hs__fill_4 FILLER_208_138 ();
 sky130_fd_sc_hs__fill_2 FILLER_208_142 ();
 sky130_fd_sc_hs__fill_1 FILLER_208_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_208_146 ();
 sky130_fd_sc_hs__fill_4 FILLER_208_154 ();
 sky130_fd_sc_hs__fill_2 FILLER_208_158 ();
 sky130_fd_sc_hs__fill_1 FILLER_208_160 ();
 sky130_fd_sc_hs__fill_2 FILLER_208_200 ();
 sky130_fd_sc_hs__fill_1 FILLER_208_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_208_225 ();
 sky130_fd_sc_hs__fill_1 FILLER_208_233 ();
 sky130_fd_sc_hs__fill_4 FILLER_208_237 ();
 sky130_fd_sc_hs__fill_2 FILLER_208_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_208_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_208_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_208_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_208_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_208_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_208_302 ();
 sky130_fd_sc_hs__fill_8 FILLER_208_310 ();
 sky130_fd_sc_hs__fill_1 FILLER_208_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_208_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_208_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_208_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_208_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_208_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_208_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_208_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_208_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_208_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_208_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_208_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_208_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_208_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_208_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_208_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_208_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_208_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_208_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_208_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_208_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_208_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_208_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_208_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_208_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_208_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_208_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_208_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_208_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_208_526 ();
 sky130_fd_sc_hs__fill_4 FILLER_208_534 ();
 sky130_fd_sc_hs__fill_2 FILLER_208_538 ();
 sky130_fd_sc_hs__fill_4 FILLER_209_0 ();
 sky130_fd_sc_hs__fill_2 FILLER_209_4 ();
 sky130_fd_sc_hs__fill_2 FILLER_209_14 ();
 sky130_fd_sc_hs__fill_1 FILLER_209_16 ();
 sky130_fd_sc_hs__fill_1 FILLER_209_25 ();
 sky130_fd_sc_hs__fill_8 FILLER_209_41 ();
 sky130_fd_sc_hs__fill_8 FILLER_209_49 ();
 sky130_fd_sc_hs__fill_1 FILLER_209_57 ();
 sky130_fd_sc_hs__fill_4 FILLER_209_59 ();
 sky130_fd_sc_hs__fill_2 FILLER_209_63 ();
 sky130_fd_sc_hs__fill_1 FILLER_209_65 ();
 sky130_fd_sc_hs__fill_8 FILLER_209_101 ();
 sky130_fd_sc_hs__fill_4 FILLER_209_109 ();
 sky130_fd_sc_hs__fill_2 FILLER_209_113 ();
 sky130_fd_sc_hs__fill_1 FILLER_209_115 ();
 sky130_fd_sc_hs__fill_2 FILLER_209_117 ();
 sky130_fd_sc_hs__fill_1 FILLER_209_119 ();
 sky130_fd_sc_hs__fill_8 FILLER_209_155 ();
 sky130_fd_sc_hs__fill_8 FILLER_209_163 ();
 sky130_fd_sc_hs__fill_2 FILLER_209_171 ();
 sky130_fd_sc_hs__fill_1 FILLER_209_173 ();
 sky130_fd_sc_hs__fill_2 FILLER_209_227 ();
 sky130_fd_sc_hs__fill_8 FILLER_209_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_209_241 ();
 sky130_fd_sc_hs__fill_1 FILLER_209_249 ();
 sky130_fd_sc_hs__fill_4 FILLER_209_276 ();
 sky130_fd_sc_hs__fill_4 FILLER_209_285 ();
 sky130_fd_sc_hs__fill_1 FILLER_209_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_209_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_209_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_209_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_209_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_209_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_209_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_209_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_209_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_209_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_209_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_209_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_209_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_209_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_209_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_209_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_209_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_209_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_209_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_209_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_209_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_209_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_209_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_209_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_209_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_209_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_209_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_209_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_209_489 ();
 sky130_fd_sc_hs__fill_1 FILLER_209_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_209_506 ();
 sky130_fd_sc_hs__fill_8 FILLER_209_514 ();
 sky130_fd_sc_hs__fill_8 FILLER_209_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_209_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_209_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_210_0 ();
 sky130_fd_sc_hs__fill_1 FILLER_210_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_210_37 ();
 sky130_fd_sc_hs__fill_8 FILLER_210_45 ();
 sky130_fd_sc_hs__fill_8 FILLER_210_53 ();
 sky130_fd_sc_hs__fill_8 FILLER_210_61 ();
 sky130_fd_sc_hs__fill_8 FILLER_210_69 ();
 sky130_fd_sc_hs__fill_8 FILLER_210_77 ();
 sky130_fd_sc_hs__fill_2 FILLER_210_85 ();
 sky130_fd_sc_hs__fill_8 FILLER_210_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_210_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_210_107 ();
 sky130_fd_sc_hs__fill_8 FILLER_210_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_210_123 ();
 sky130_fd_sc_hs__fill_8 FILLER_210_131 ();
 sky130_fd_sc_hs__fill_4 FILLER_210_139 ();
 sky130_fd_sc_hs__fill_2 FILLER_210_143 ();
 sky130_fd_sc_hs__fill_8 FILLER_210_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_210_154 ();
 sky130_fd_sc_hs__fill_1 FILLER_210_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_210_184 ();
 sky130_fd_sc_hs__fill_8 FILLER_210_192 ();
 sky130_fd_sc_hs__fill_2 FILLER_210_200 ();
 sky130_fd_sc_hs__fill_1 FILLER_210_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_210_225 ();
 sky130_fd_sc_hs__fill_4 FILLER_210_233 ();
 sky130_fd_sc_hs__fill_2 FILLER_210_237 ();
 sky130_fd_sc_hs__fill_1 FILLER_210_239 ();
 sky130_fd_sc_hs__fill_8 FILLER_210_262 ();
 sky130_fd_sc_hs__fill_4 FILLER_210_270 ();
 sky130_fd_sc_hs__fill_1 FILLER_210_274 ();
 sky130_fd_sc_hs__fill_4 FILLER_210_312 ();
 sky130_fd_sc_hs__fill_2 FILLER_210_316 ();
 sky130_fd_sc_hs__fill_1 FILLER_210_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_210_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_210_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_210_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_210_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_210_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_210_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_210_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_210_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_210_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_210_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_210_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_210_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_210_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_210_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_210_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_210_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_210_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_210_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_210_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_210_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_210_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_210_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_210_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_210_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_210_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_210_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_210_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_210_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_210_526 ();
 sky130_fd_sc_hs__fill_4 FILLER_210_534 ();
 sky130_fd_sc_hs__fill_2 FILLER_210_538 ();
 sky130_fd_sc_hs__fill_8 FILLER_211_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_211_8 ();
 sky130_fd_sc_hs__fill_4 FILLER_211_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_211_25 ();
 sky130_fd_sc_hs__fill_2 FILLER_211_29 ();
 sky130_fd_sc_hs__fill_4 FILLER_211_34 ();
 sky130_fd_sc_hs__fill_2 FILLER_211_38 ();
 sky130_fd_sc_hs__fill_1 FILLER_211_40 ();
 sky130_fd_sc_hs__fill_8 FILLER_211_50 ();
 sky130_fd_sc_hs__fill_2 FILLER_211_59 ();
 sky130_fd_sc_hs__fill_1 FILLER_211_61 ();
 sky130_fd_sc_hs__fill_8 FILLER_211_79 ();
 sky130_fd_sc_hs__fill_8 FILLER_211_87 ();
 sky130_fd_sc_hs__fill_8 FILLER_211_95 ();
 sky130_fd_sc_hs__fill_8 FILLER_211_103 ();
 sky130_fd_sc_hs__fill_4 FILLER_211_111 ();
 sky130_fd_sc_hs__fill_1 FILLER_211_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_211_117 ();
 sky130_fd_sc_hs__fill_4 FILLER_211_125 ();
 sky130_fd_sc_hs__fill_2 FILLER_211_129 ();
 sky130_fd_sc_hs__fill_8 FILLER_211_166 ();
 sky130_fd_sc_hs__fill_8 FILLER_211_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_211_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_211_191 ();
 sky130_fd_sc_hs__fill_4 FILLER_211_199 ();
 sky130_fd_sc_hs__fill_2 FILLER_211_203 ();
 sky130_fd_sc_hs__fill_1 FILLER_211_205 ();
 sky130_fd_sc_hs__fill_8 FILLER_211_219 ();
 sky130_fd_sc_hs__fill_4 FILLER_211_227 ();
 sky130_fd_sc_hs__fill_1 FILLER_211_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_211_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_211_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_211_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_211_268 ();
 sky130_fd_sc_hs__fill_8 FILLER_211_276 ();
 sky130_fd_sc_hs__fill_4 FILLER_211_284 ();
 sky130_fd_sc_hs__fill_2 FILLER_211_288 ();
 sky130_fd_sc_hs__fill_8 FILLER_211_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_211_317 ();
 sky130_fd_sc_hs__fill_8 FILLER_211_325 ();
 sky130_fd_sc_hs__fill_8 FILLER_211_333 ();
 sky130_fd_sc_hs__fill_4 FILLER_211_341 ();
 sky130_fd_sc_hs__fill_2 FILLER_211_345 ();
 sky130_fd_sc_hs__fill_1 FILLER_211_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_211_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_211_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_211_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_211_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_211_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_211_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_211_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_211_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_211_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_211_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_211_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_211_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_211_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_211_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_211_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_211_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_211_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_211_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_211_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_211_489 ();
 sky130_fd_sc_hs__fill_1 FILLER_211_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_211_506 ();
 sky130_fd_sc_hs__fill_8 FILLER_211_514 ();
 sky130_fd_sc_hs__fill_8 FILLER_211_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_211_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_211_539 ();
 sky130_fd_sc_hs__fill_2 FILLER_212_8 ();
 sky130_fd_sc_hs__fill_1 FILLER_212_10 ();
 sky130_fd_sc_hs__fill_2 FILLER_212_30 ();
 sky130_fd_sc_hs__fill_2 FILLER_212_40 ();
 sky130_fd_sc_hs__fill_4 FILLER_212_74 ();
 sky130_fd_sc_hs__fill_2 FILLER_212_78 ();
 sky130_fd_sc_hs__fill_4 FILLER_212_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_212_88 ();
 sky130_fd_sc_hs__fill_4 FILLER_212_96 ();
 sky130_fd_sc_hs__fill_2 FILLER_212_100 ();
 sky130_fd_sc_hs__fill_1 FILLER_212_102 ();
 sky130_fd_sc_hs__fill_4 FILLER_212_138 ();
 sky130_fd_sc_hs__fill_2 FILLER_212_142 ();
 sky130_fd_sc_hs__fill_1 FILLER_212_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_212_146 ();
 sky130_fd_sc_hs__fill_4 FILLER_212_154 ();
 sky130_fd_sc_hs__fill_2 FILLER_212_158 ();
 sky130_fd_sc_hs__fill_1 FILLER_212_160 ();
 sky130_fd_sc_hs__fill_8 FILLER_212_182 ();
 sky130_fd_sc_hs__fill_8 FILLER_212_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_212_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_212_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_212_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_212_236 ();
 sky130_fd_sc_hs__fill_1 FILLER_212_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_212_253 ();
 sky130_fd_sc_hs__fill_8 FILLER_212_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_212_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_212_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_212_286 ();
 sky130_fd_sc_hs__fill_4 FILLER_212_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_212_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_212_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_212_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_212_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_212_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_212_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_212_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_212_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_212_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_212_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_212_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_212_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_212_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_212_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_212_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_212_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_212_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_212_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_212_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_212_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_212_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_212_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_212_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_212_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_212_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_212_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_212_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_212_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_212_526 ();
 sky130_fd_sc_hs__fill_4 FILLER_212_534 ();
 sky130_fd_sc_hs__fill_2 FILLER_212_538 ();
 sky130_fd_sc_hs__fill_8 FILLER_213_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_213_16 ();
 sky130_fd_sc_hs__fill_2 FILLER_213_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_213_26 ();
 sky130_fd_sc_hs__fill_8 FILLER_213_38 ();
 sky130_fd_sc_hs__fill_2 FILLER_213_46 ();
 sky130_fd_sc_hs__fill_1 FILLER_213_48 ();
 sky130_fd_sc_hs__fill_4 FILLER_213_52 ();
 sky130_fd_sc_hs__fill_2 FILLER_213_56 ();
 sky130_fd_sc_hs__fill_4 FILLER_213_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_213_75 ();
 sky130_fd_sc_hs__fill_1 FILLER_213_83 ();
 sky130_fd_sc_hs__fill_4 FILLER_213_105 ();
 sky130_fd_sc_hs__fill_1 FILLER_213_109 ();
 sky130_fd_sc_hs__fill_1 FILLER_213_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_213_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_213_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_213_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_213_141 ();
 sky130_fd_sc_hs__fill_4 FILLER_213_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_213_175 ();
 sky130_fd_sc_hs__fill_2 FILLER_213_183 ();
 sky130_fd_sc_hs__fill_1 FILLER_213_185 ();
 sky130_fd_sc_hs__fill_4 FILLER_213_195 ();
 sky130_fd_sc_hs__fill_8 FILLER_213_220 ();
 sky130_fd_sc_hs__fill_4 FILLER_213_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_213_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_213_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_213_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_213_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_213_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_213_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_213_281 ();
 sky130_fd_sc_hs__fill_1 FILLER_213_289 ();
 sky130_fd_sc_hs__fill_8 FILLER_213_291 ();
 sky130_fd_sc_hs__fill_1 FILLER_213_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_213_305 ();
 sky130_fd_sc_hs__fill_8 FILLER_213_313 ();
 sky130_fd_sc_hs__fill_8 FILLER_213_321 ();
 sky130_fd_sc_hs__fill_8 FILLER_213_329 ();
 sky130_fd_sc_hs__fill_8 FILLER_213_337 ();
 sky130_fd_sc_hs__fill_2 FILLER_213_345 ();
 sky130_fd_sc_hs__fill_1 FILLER_213_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_213_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_213_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_213_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_213_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_213_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_213_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_213_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_213_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_213_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_213_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_213_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_213_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_213_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_213_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_213_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_213_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_213_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_213_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_213_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_213_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_213_500 ();
 sky130_fd_sc_hs__fill_1 FILLER_213_508 ();
 sky130_fd_sc_hs__fill_8 FILLER_213_512 ();
 sky130_fd_sc_hs__fill_2 FILLER_213_520 ();
 sky130_fd_sc_hs__fill_4 FILLER_213_523 ();
 sky130_fd_sc_hs__fill_4 FILLER_213_535 ();
 sky130_fd_sc_hs__fill_1 FILLER_213_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_214_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_214_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_214_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_214_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_214_28 ();
 sky130_fd_sc_hs__fill_4 FILLER_214_35 ();
 sky130_fd_sc_hs__fill_1 FILLER_214_39 ();
 sky130_fd_sc_hs__fill_8 FILLER_214_57 ();
 sky130_fd_sc_hs__fill_8 FILLER_214_65 ();
 sky130_fd_sc_hs__fill_2 FILLER_214_73 ();
 sky130_fd_sc_hs__fill_8 FILLER_214_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_214_96 ();
 sky130_fd_sc_hs__fill_4 FILLER_214_104 ();
 sky130_fd_sc_hs__fill_2 FILLER_214_108 ();
 sky130_fd_sc_hs__fill_2 FILLER_214_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_214_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_214_165 ();
 sky130_fd_sc_hs__fill_8 FILLER_214_173 ();
 sky130_fd_sc_hs__fill_1 FILLER_214_181 ();
 sky130_fd_sc_hs__fill_8 FILLER_214_204 ();
 sky130_fd_sc_hs__fill_4 FILLER_214_212 ();
 sky130_fd_sc_hs__fill_1 FILLER_214_216 ();
 sky130_fd_sc_hs__fill_2 FILLER_214_259 ();
 sky130_fd_sc_hs__fill_8 FILLER_214_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_214_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_214_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_214_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_214_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_214_302 ();
 sky130_fd_sc_hs__fill_8 FILLER_214_310 ();
 sky130_fd_sc_hs__fill_1 FILLER_214_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_214_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_214_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_214_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_214_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_214_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_214_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_214_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_214_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_214_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_214_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_214_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_214_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_214_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_214_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_214_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_214_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_214_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_214_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_214_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_214_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_214_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_214_476 ();
 sky130_fd_sc_hs__fill_2 FILLER_214_484 ();
 sky130_fd_sc_hs__fill_4 FILLER_214_494 ();
 sky130_fd_sc_hs__fill_1 FILLER_214_498 ();
 sky130_fd_sc_hs__fill_8 FILLER_214_514 ();
 sky130_fd_sc_hs__fill_8 FILLER_214_522 ();
 sky130_fd_sc_hs__fill_8 FILLER_214_530 ();
 sky130_fd_sc_hs__fill_2 FILLER_214_538 ();
 sky130_fd_sc_hs__fill_4 FILLER_215_8 ();
 sky130_fd_sc_hs__fill_1 FILLER_215_12 ();
 sky130_fd_sc_hs__fill_2 FILLER_215_26 ();
 sky130_fd_sc_hs__fill_4 FILLER_215_35 ();
 sky130_fd_sc_hs__fill_1 FILLER_215_39 ();
 sky130_fd_sc_hs__fill_4 FILLER_215_53 ();
 sky130_fd_sc_hs__fill_1 FILLER_215_57 ();
 sky130_fd_sc_hs__fill_8 FILLER_215_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_215_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_215_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_215_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_215_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_215_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_215_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_215_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_215_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_215_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_215_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_215_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_215_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_215_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_215_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_215_173 ();
 sky130_fd_sc_hs__fill_2 FILLER_215_175 ();
 sky130_fd_sc_hs__fill_1 FILLER_215_177 ();
 sky130_fd_sc_hs__fill_8 FILLER_215_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_215_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_215_215 ();
 sky130_fd_sc_hs__fill_4 FILLER_215_223 ();
 sky130_fd_sc_hs__fill_2 FILLER_215_227 ();
 sky130_fd_sc_hs__fill_2 FILLER_215_242 ();
 sky130_fd_sc_hs__fill_1 FILLER_215_244 ();
 sky130_fd_sc_hs__fill_2 FILLER_215_251 ();
 sky130_fd_sc_hs__fill_1 FILLER_215_253 ();
 sky130_fd_sc_hs__fill_2 FILLER_215_267 ();
 sky130_fd_sc_hs__fill_8 FILLER_215_279 ();
 sky130_fd_sc_hs__fill_2 FILLER_215_287 ();
 sky130_fd_sc_hs__fill_1 FILLER_215_289 ();
 sky130_fd_sc_hs__fill_4 FILLER_215_291 ();
 sky130_fd_sc_hs__fill_1 FILLER_215_295 ();
 sky130_fd_sc_hs__fill_8 FILLER_215_301 ();
 sky130_fd_sc_hs__fill_8 FILLER_215_309 ();
 sky130_fd_sc_hs__fill_8 FILLER_215_317 ();
 sky130_fd_sc_hs__fill_8 FILLER_215_325 ();
 sky130_fd_sc_hs__fill_8 FILLER_215_333 ();
 sky130_fd_sc_hs__fill_4 FILLER_215_341 ();
 sky130_fd_sc_hs__fill_2 FILLER_215_345 ();
 sky130_fd_sc_hs__fill_1 FILLER_215_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_215_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_215_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_215_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_215_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_215_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_215_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_215_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_215_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_215_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_215_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_215_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_215_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_215_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_215_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_215_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_215_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_215_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_215_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_215_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_215_489 ();
 sky130_fd_sc_hs__fill_1 FILLER_215_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_215_506 ();
 sky130_fd_sc_hs__fill_8 FILLER_215_514 ();
 sky130_fd_sc_hs__fill_8 FILLER_215_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_215_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_215_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_216_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_216_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_216_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_216_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_216_28 ();
 sky130_fd_sc_hs__fill_4 FILLER_216_30 ();
 sky130_fd_sc_hs__fill_2 FILLER_216_34 ();
 sky130_fd_sc_hs__fill_8 FILLER_216_41 ();
 sky130_fd_sc_hs__fill_8 FILLER_216_49 ();
 sky130_fd_sc_hs__fill_8 FILLER_216_57 ();
 sky130_fd_sc_hs__fill_8 FILLER_216_65 ();
 sky130_fd_sc_hs__fill_8 FILLER_216_73 ();
 sky130_fd_sc_hs__fill_4 FILLER_216_81 ();
 sky130_fd_sc_hs__fill_2 FILLER_216_85 ();
 sky130_fd_sc_hs__fill_4 FILLER_216_88 ();
 sky130_fd_sc_hs__fill_2 FILLER_216_92 ();
 sky130_fd_sc_hs__fill_4 FILLER_216_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_216_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_216_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_216_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_216_170 ();
 sky130_fd_sc_hs__fill_4 FILLER_216_178 ();
 sky130_fd_sc_hs__fill_2 FILLER_216_182 ();
 sky130_fd_sc_hs__fill_1 FILLER_216_184 ();
 sky130_fd_sc_hs__fill_4 FILLER_216_204 ();
 sky130_fd_sc_hs__fill_2 FILLER_216_208 ();
 sky130_fd_sc_hs__fill_8 FILLER_216_213 ();
 sky130_fd_sc_hs__fill_8 FILLER_216_221 ();
 sky130_fd_sc_hs__fill_8 FILLER_216_229 ();
 sky130_fd_sc_hs__fill_2 FILLER_216_237 ();
 sky130_fd_sc_hs__fill_1 FILLER_216_239 ();
 sky130_fd_sc_hs__fill_8 FILLER_216_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_216_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_216_278 ();
 sky130_fd_sc_hs__fill_4 FILLER_216_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_216_311 ();
 sky130_fd_sc_hs__fill_8 FILLER_216_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_216_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_216_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_216_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_216_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_216_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_216_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_216_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_216_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_216_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_216_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_216_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_216_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_216_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_216_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_216_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_216_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_216_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_216_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_216_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_216_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_216_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_216_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_216_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_216_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_216_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_216_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_216_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_216_526 ();
 sky130_fd_sc_hs__fill_4 FILLER_216_534 ();
 sky130_fd_sc_hs__fill_2 FILLER_216_538 ();
 sky130_fd_sc_hs__fill_8 FILLER_217_0 ();
 sky130_fd_sc_hs__fill_4 FILLER_217_8 ();
 sky130_fd_sc_hs__fill_2 FILLER_217_12 ();
 sky130_fd_sc_hs__fill_8 FILLER_217_22 ();
 sky130_fd_sc_hs__fill_2 FILLER_217_30 ();
 sky130_fd_sc_hs__fill_2 FILLER_217_44 ();
 sky130_fd_sc_hs__fill_8 FILLER_217_59 ();
 sky130_fd_sc_hs__fill_4 FILLER_217_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_217_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_217_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_217_104 ();
 sky130_fd_sc_hs__fill_4 FILLER_217_112 ();
 sky130_fd_sc_hs__fill_4 FILLER_217_117 ();
 sky130_fd_sc_hs__fill_1 FILLER_217_121 ();
 sky130_fd_sc_hs__fill_8 FILLER_217_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_217_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_217_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_217_175 ();
 sky130_fd_sc_hs__fill_4 FILLER_217_183 ();
 sky130_fd_sc_hs__fill_1 FILLER_217_187 ();
 sky130_fd_sc_hs__fill_8 FILLER_217_193 ();
 sky130_fd_sc_hs__fill_4 FILLER_217_201 ();
 sky130_fd_sc_hs__fill_2 FILLER_217_205 ();
 sky130_fd_sc_hs__fill_1 FILLER_217_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_217_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_217_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_217_254 ();
 sky130_fd_sc_hs__fill_8 FILLER_217_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_217_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_217_278 ();
 sky130_fd_sc_hs__fill_4 FILLER_217_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_217_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_217_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_217_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_217_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_217_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_217_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_217_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_217_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_217_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_217_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_217_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_217_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_217_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_217_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_217_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_217_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_217_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_217_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_217_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_217_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_217_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_217_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_217_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_217_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_217_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_217_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_217_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_217_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_217_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_217_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_217_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_217_521 ();
 sky130_fd_sc_hs__fill_2 FILLER_217_523 ();
 sky130_fd_sc_hs__fill_4 FILLER_217_533 ();
 sky130_fd_sc_hs__fill_2 FILLER_217_537 ();
 sky130_fd_sc_hs__fill_1 FILLER_217_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_218_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_218_8 ();
 sky130_fd_sc_hs__fill_4 FILLER_218_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_218_28 ();
 sky130_fd_sc_hs__fill_4 FILLER_218_30 ();
 sky130_fd_sc_hs__fill_2 FILLER_218_34 ();
 sky130_fd_sc_hs__fill_8 FILLER_218_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_218_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_218_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_218_96 ();
 sky130_fd_sc_hs__fill_8 FILLER_218_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_218_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_218_120 ();
 sky130_fd_sc_hs__fill_8 FILLER_218_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_218_136 ();
 sky130_fd_sc_hs__fill_1 FILLER_218_144 ();
 sky130_fd_sc_hs__fill_8 FILLER_218_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_218_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_218_162 ();
 sky130_fd_sc_hs__fill_4 FILLER_218_170 ();
 sky130_fd_sc_hs__fill_4 FILLER_218_199 ();
 sky130_fd_sc_hs__fill_2 FILLER_218_204 ();
 sky130_fd_sc_hs__fill_1 FILLER_218_206 ();
 sky130_fd_sc_hs__fill_8 FILLER_218_214 ();
 sky130_fd_sc_hs__fill_8 FILLER_218_222 ();
 sky130_fd_sc_hs__fill_8 FILLER_218_230 ();
 sky130_fd_sc_hs__fill_2 FILLER_218_238 ();
 sky130_fd_sc_hs__fill_8 FILLER_218_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_218_270 ();
 sky130_fd_sc_hs__fill_2 FILLER_218_278 ();
 sky130_fd_sc_hs__fill_1 FILLER_218_280 ();
 sky130_fd_sc_hs__fill_2 FILLER_218_293 ();
 sky130_fd_sc_hs__fill_1 FILLER_218_295 ();
 sky130_fd_sc_hs__fill_8 FILLER_218_309 ();
 sky130_fd_sc_hs__fill_2 FILLER_218_317 ();
 sky130_fd_sc_hs__fill_8 FILLER_218_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_218_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_218_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_218_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_218_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_218_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_218_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_218_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_218_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_218_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_218_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_218_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_218_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_218_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_218_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_218_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_218_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_218_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_218_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_218_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_218_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_218_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_218_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_218_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_218_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_218_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_218_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_218_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_218_526 ();
 sky130_fd_sc_hs__fill_4 FILLER_218_534 ();
 sky130_fd_sc_hs__fill_2 FILLER_218_538 ();
 sky130_fd_sc_hs__fill_8 FILLER_219_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_219_8 ();
 sky130_fd_sc_hs__fill_4 FILLER_219_16 ();
 sky130_fd_sc_hs__fill_2 FILLER_219_20 ();
 sky130_fd_sc_hs__fill_8 FILLER_219_30 ();
 sky130_fd_sc_hs__fill_4 FILLER_219_38 ();
 sky130_fd_sc_hs__fill_1 FILLER_219_42 ();
 sky130_fd_sc_hs__fill_8 FILLER_219_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_219_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_219_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_219_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_219_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_219_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_219_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_219_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_219_117 ();
 sky130_fd_sc_hs__fill_4 FILLER_219_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_219_164 ();
 sky130_fd_sc_hs__fill_2 FILLER_219_172 ();
 sky130_fd_sc_hs__fill_2 FILLER_219_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_219_198 ();
 sky130_fd_sc_hs__fill_4 FILLER_219_206 ();
 sky130_fd_sc_hs__fill_1 FILLER_219_210 ();
 sky130_fd_sc_hs__fill_8 FILLER_219_233 ();
 sky130_fd_sc_hs__fill_4 FILLER_219_241 ();
 sky130_fd_sc_hs__fill_2 FILLER_219_245 ();
 sky130_fd_sc_hs__fill_1 FILLER_219_247 ();
 sky130_fd_sc_hs__fill_1 FILLER_219_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_219_305 ();
 sky130_fd_sc_hs__fill_8 FILLER_219_313 ();
 sky130_fd_sc_hs__fill_8 FILLER_219_321 ();
 sky130_fd_sc_hs__fill_8 FILLER_219_329 ();
 sky130_fd_sc_hs__fill_8 FILLER_219_337 ();
 sky130_fd_sc_hs__fill_2 FILLER_219_345 ();
 sky130_fd_sc_hs__fill_1 FILLER_219_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_219_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_219_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_219_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_219_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_219_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_219_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_219_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_219_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_219_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_219_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_219_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_219_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_219_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_219_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_219_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_219_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_219_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_219_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_219_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_219_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_219_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_219_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_219_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_219_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_219_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_219_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_219_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_220_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_220_28 ();
 sky130_fd_sc_hs__fill_4 FILLER_220_30 ();
 sky130_fd_sc_hs__fill_2 FILLER_220_34 ();
 sky130_fd_sc_hs__fill_1 FILLER_220_36 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_64 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_72 ();
 sky130_fd_sc_hs__fill_4 FILLER_220_80 ();
 sky130_fd_sc_hs__fill_2 FILLER_220_84 ();
 sky130_fd_sc_hs__fill_1 FILLER_220_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_96 ();
 sky130_fd_sc_hs__fill_4 FILLER_220_104 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_113 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_121 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_129 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_137 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_178 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_186 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_194 ();
 sky130_fd_sc_hs__fill_1 FILLER_220_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_236 ();
 sky130_fd_sc_hs__fill_4 FILLER_220_244 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_270 ();
 sky130_fd_sc_hs__fill_4 FILLER_220_278 ();
 sky130_fd_sc_hs__fill_1 FILLER_220_282 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_304 ();
 sky130_fd_sc_hs__fill_4 FILLER_220_312 ();
 sky130_fd_sc_hs__fill_2 FILLER_220_316 ();
 sky130_fd_sc_hs__fill_1 FILLER_220_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_220_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_220_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_220_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_220_526 ();
 sky130_fd_sc_hs__fill_4 FILLER_220_534 ();
 sky130_fd_sc_hs__fill_2 FILLER_220_538 ();
 sky130_fd_sc_hs__fill_8 FILLER_221_0 ();
 sky130_fd_sc_hs__fill_4 FILLER_221_8 ();
 sky130_fd_sc_hs__fill_2 FILLER_221_12 ();
 sky130_fd_sc_hs__fill_8 FILLER_221_22 ();
 sky130_fd_sc_hs__fill_8 FILLER_221_30 ();
 sky130_fd_sc_hs__fill_2 FILLER_221_38 ();
 sky130_fd_sc_hs__fill_1 FILLER_221_40 ();
 sky130_fd_sc_hs__fill_2 FILLER_221_56 ();
 sky130_fd_sc_hs__fill_8 FILLER_221_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_221_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_221_75 ();
 sky130_fd_sc_hs__fill_2 FILLER_221_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_221_98 ();
 sky130_fd_sc_hs__fill_2 FILLER_221_106 ();
 sky130_fd_sc_hs__fill_1 FILLER_221_108 ();
 sky130_fd_sc_hs__fill_4 FILLER_221_112 ();
 sky130_fd_sc_hs__fill_8 FILLER_221_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_221_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_221_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_221_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_221_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_221_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_221_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_221_173 ();
 sky130_fd_sc_hs__fill_2 FILLER_221_175 ();
 sky130_fd_sc_hs__fill_1 FILLER_221_177 ();
 sky130_fd_sc_hs__fill_8 FILLER_221_199 ();
 sky130_fd_sc_hs__fill_4 FILLER_221_207 ();
 sky130_fd_sc_hs__fill_4 FILLER_221_246 ();
 sky130_fd_sc_hs__fill_8 FILLER_221_266 ();
 sky130_fd_sc_hs__fill_8 FILLER_221_274 ();
 sky130_fd_sc_hs__fill_8 FILLER_221_282 ();
 sky130_fd_sc_hs__fill_8 FILLER_221_309 ();
 sky130_fd_sc_hs__fill_8 FILLER_221_317 ();
 sky130_fd_sc_hs__fill_8 FILLER_221_325 ();
 sky130_fd_sc_hs__fill_8 FILLER_221_333 ();
 sky130_fd_sc_hs__fill_4 FILLER_221_341 ();
 sky130_fd_sc_hs__fill_2 FILLER_221_345 ();
 sky130_fd_sc_hs__fill_1 FILLER_221_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_221_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_221_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_221_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_221_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_221_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_221_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_221_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_221_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_221_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_221_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_221_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_221_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_221_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_221_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_221_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_221_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_221_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_221_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_221_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_221_489 ();
 sky130_fd_sc_hs__fill_1 FILLER_221_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_221_506 ();
 sky130_fd_sc_hs__fill_8 FILLER_221_514 ();
 sky130_fd_sc_hs__fill_8 FILLER_221_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_221_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_221_539 ();
 sky130_fd_sc_hs__fill_4 FILLER_222_0 ();
 sky130_fd_sc_hs__fill_2 FILLER_222_4 ();
 sky130_fd_sc_hs__fill_1 FILLER_222_6 ();
 sky130_fd_sc_hs__fill_8 FILLER_222_15 ();
 sky130_fd_sc_hs__fill_4 FILLER_222_23 ();
 sky130_fd_sc_hs__fill_2 FILLER_222_27 ();
 sky130_fd_sc_hs__fill_8 FILLER_222_30 ();
 sky130_fd_sc_hs__fill_4 FILLER_222_38 ();
 sky130_fd_sc_hs__fill_2 FILLER_222_42 ();
 sky130_fd_sc_hs__fill_8 FILLER_222_55 ();
 sky130_fd_sc_hs__fill_8 FILLER_222_63 ();
 sky130_fd_sc_hs__fill_8 FILLER_222_71 ();
 sky130_fd_sc_hs__fill_2 FILLER_222_79 ();
 sky130_fd_sc_hs__fill_1 FILLER_222_81 ();
 sky130_fd_sc_hs__fill_8 FILLER_222_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_222_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_222_133 ();
 sky130_fd_sc_hs__fill_4 FILLER_222_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_222_167 ();
 sky130_fd_sc_hs__fill_8 FILLER_222_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_222_183 ();
 sky130_fd_sc_hs__fill_4 FILLER_222_191 ();
 sky130_fd_sc_hs__fill_1 FILLER_222_195 ();
 sky130_fd_sc_hs__fill_2 FILLER_222_201 ();
 sky130_fd_sc_hs__fill_1 FILLER_222_204 ();
 sky130_fd_sc_hs__fill_2 FILLER_222_226 ();
 sky130_fd_sc_hs__fill_1 FILLER_222_228 ();
 sky130_fd_sc_hs__fill_8 FILLER_222_249 ();
 sky130_fd_sc_hs__fill_4 FILLER_222_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_222_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_222_270 ();
 sky130_fd_sc_hs__fill_1 FILLER_222_278 ();
 sky130_fd_sc_hs__fill_2 FILLER_222_292 ();
 sky130_fd_sc_hs__fill_1 FILLER_222_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_222_307 ();
 sky130_fd_sc_hs__fill_4 FILLER_222_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_222_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_222_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_222_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_222_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_222_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_222_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_222_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_222_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_222_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_222_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_222_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_222_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_222_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_222_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_222_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_222_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_222_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_222_444 ();
 sky130_fd_sc_hs__fill_8 FILLER_222_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_222_460 ();
 sky130_fd_sc_hs__fill_8 FILLER_222_468 ();
 sky130_fd_sc_hs__fill_8 FILLER_222_476 ();
 sky130_fd_sc_hs__fill_8 FILLER_222_484 ();
 sky130_fd_sc_hs__fill_1 FILLER_222_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_222_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_222_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_222_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_222_526 ();
 sky130_fd_sc_hs__fill_4 FILLER_222_534 ();
 sky130_fd_sc_hs__fill_2 FILLER_222_538 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_0 ();
 sky130_fd_sc_hs__fill_4 FILLER_223_8 ();
 sky130_fd_sc_hs__fill_1 FILLER_223_12 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_21 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_29 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_37 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_45 ();
 sky130_fd_sc_hs__fill_4 FILLER_223_53 ();
 sky130_fd_sc_hs__fill_1 FILLER_223_57 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_59 ();
 sky130_fd_sc_hs__fill_4 FILLER_223_67 ();
 sky130_fd_sc_hs__fill_2 FILLER_223_71 ();
 sky130_fd_sc_hs__fill_1 FILLER_223_73 ();
 sky130_fd_sc_hs__fill_4 FILLER_223_91 ();
 sky130_fd_sc_hs__fill_1 FILLER_223_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_149 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_157 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_165 ();
 sky130_fd_sc_hs__fill_1 FILLER_223_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_191 ();
 sky130_fd_sc_hs__fill_4 FILLER_223_199 ();
 sky130_fd_sc_hs__fill_1 FILLER_223_203 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_221 ();
 sky130_fd_sc_hs__fill_2 FILLER_223_229 ();
 sky130_fd_sc_hs__fill_1 FILLER_223_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_257 ();
 sky130_fd_sc_hs__fill_4 FILLER_223_265 ();
 sky130_fd_sc_hs__fill_2 FILLER_223_269 ();
 sky130_fd_sc_hs__fill_1 FILLER_223_271 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_223_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_381 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_389 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_397 ();
 sky130_fd_sc_hs__fill_1 FILLER_223_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_447 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_455 ();
 sky130_fd_sc_hs__fill_1 FILLER_223_463 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_489 ();
 sky130_fd_sc_hs__fill_1 FILLER_223_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_506 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_514 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_223_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_223_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_224_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_224_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_38 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_54 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_62 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_70 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_78 ();
 sky130_fd_sc_hs__fill_1 FILLER_224_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_88 ();
 sky130_fd_sc_hs__fill_4 FILLER_224_96 ();
 sky130_fd_sc_hs__fill_2 FILLER_224_100 ();
 sky130_fd_sc_hs__fill_1 FILLER_224_102 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_124 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_132 ();
 sky130_fd_sc_hs__fill_4 FILLER_224_140 ();
 sky130_fd_sc_hs__fill_1 FILLER_224_144 ();
 sky130_fd_sc_hs__fill_2 FILLER_224_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_169 ();
 sky130_fd_sc_hs__fill_4 FILLER_224_198 ();
 sky130_fd_sc_hs__fill_1 FILLER_224_202 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_212 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_228 ();
 sky130_fd_sc_hs__fill_4 FILLER_224_236 ();
 sky130_fd_sc_hs__fill_1 FILLER_224_240 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_248 ();
 sky130_fd_sc_hs__fill_4 FILLER_224_256 ();
 sky130_fd_sc_hs__fill_1 FILLER_224_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_262 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_270 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_278 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_286 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_294 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_302 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_310 ();
 sky130_fd_sc_hs__fill_1 FILLER_224_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_224_376 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_378 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_386 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_394 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_402 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_410 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_418 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_426 ();
 sky130_fd_sc_hs__fill_1 FILLER_224_434 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_444 ();
 sky130_fd_sc_hs__fill_4 FILLER_224_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_458 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_466 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_474 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_482 ();
 sky130_fd_sc_hs__fill_2 FILLER_224_490 ();
 sky130_fd_sc_hs__fill_1 FILLER_224_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_224_526 ();
 sky130_fd_sc_hs__fill_4 FILLER_224_534 ();
 sky130_fd_sc_hs__fill_2 FILLER_224_538 ();
 sky130_fd_sc_hs__fill_8 FILLER_225_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_225_8 ();
 sky130_fd_sc_hs__fill_4 FILLER_225_16 ();
 sky130_fd_sc_hs__fill_1 FILLER_225_20 ();
 sky130_fd_sc_hs__fill_8 FILLER_225_29 ();
 sky130_fd_sc_hs__fill_8 FILLER_225_37 ();
 sky130_fd_sc_hs__fill_4 FILLER_225_45 ();
 sky130_fd_sc_hs__fill_1 FILLER_225_49 ();
 sky130_fd_sc_hs__fill_1 FILLER_225_57 ();
 sky130_fd_sc_hs__fill_8 FILLER_225_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_225_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_225_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_225_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_225_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_225_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_225_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_225_115 ();
 sky130_fd_sc_hs__fill_8 FILLER_225_117 ();
 sky130_fd_sc_hs__fill_4 FILLER_225_125 ();
 sky130_fd_sc_hs__fill_2 FILLER_225_129 ();
 sky130_fd_sc_hs__fill_1 FILLER_225_152 ();
 sky130_fd_sc_hs__fill_4 FILLER_225_175 ();
 sky130_fd_sc_hs__fill_1 FILLER_225_179 ();
 sky130_fd_sc_hs__fill_8 FILLER_225_201 ();
 sky130_fd_sc_hs__fill_8 FILLER_225_209 ();
 sky130_fd_sc_hs__fill_8 FILLER_225_217 ();
 sky130_fd_sc_hs__fill_4 FILLER_225_225 ();
 sky130_fd_sc_hs__fill_2 FILLER_225_229 ();
 sky130_fd_sc_hs__fill_1 FILLER_225_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_225_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_225_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_225_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_225_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_225_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_225_273 ();
 sky130_fd_sc_hs__fill_8 FILLER_225_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_225_299 ();
 sky130_fd_sc_hs__fill_8 FILLER_225_307 ();
 sky130_fd_sc_hs__fill_8 FILLER_225_315 ();
 sky130_fd_sc_hs__fill_8 FILLER_225_323 ();
 sky130_fd_sc_hs__fill_8 FILLER_225_331 ();
 sky130_fd_sc_hs__fill_8 FILLER_225_339 ();
 sky130_fd_sc_hs__fill_1 FILLER_225_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_225_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_225_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_225_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_225_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_225_383 ();
 sky130_fd_sc_hs__fill_8 FILLER_225_391 ();
 sky130_fd_sc_hs__fill_4 FILLER_225_399 ();
 sky130_fd_sc_hs__fill_2 FILLER_225_403 ();
 sky130_fd_sc_hs__fill_1 FILLER_225_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_225_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_225_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_225_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_225_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_225_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_225_447 ();
 sky130_fd_sc_hs__fill_1 FILLER_225_455 ();
 sky130_fd_sc_hs__fill_4 FILLER_225_458 ();
 sky130_fd_sc_hs__fill_2 FILLER_225_462 ();
 sky130_fd_sc_hs__fill_8 FILLER_225_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_225_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_225_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_225_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_225_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_225_505 ();
 sky130_fd_sc_hs__fill_1 FILLER_225_513 ();
 sky130_fd_sc_hs__fill_8 FILLER_225_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_225_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_225_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_226_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_226_8 ();
 sky130_fd_sc_hs__fill_1 FILLER_226_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_226_25 ();
 sky130_fd_sc_hs__fill_8 FILLER_226_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_226_38 ();
 sky130_fd_sc_hs__fill_4 FILLER_226_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_226_57 ();
 sky130_fd_sc_hs__fill_8 FILLER_226_65 ();
 sky130_fd_sc_hs__fill_8 FILLER_226_73 ();
 sky130_fd_sc_hs__fill_4 FILLER_226_81 ();
 sky130_fd_sc_hs__fill_2 FILLER_226_85 ();
 sky130_fd_sc_hs__fill_2 FILLER_226_88 ();
 sky130_fd_sc_hs__fill_1 FILLER_226_90 ();
 sky130_fd_sc_hs__fill_8 FILLER_226_113 ();
 sky130_fd_sc_hs__fill_8 FILLER_226_121 ();
 sky130_fd_sc_hs__fill_8 FILLER_226_129 ();
 sky130_fd_sc_hs__fill_8 FILLER_226_137 ();
 sky130_fd_sc_hs__fill_8 FILLER_226_146 ();
 sky130_fd_sc_hs__fill_4 FILLER_226_175 ();
 sky130_fd_sc_hs__fill_1 FILLER_226_179 ();
 sky130_fd_sc_hs__fill_2 FILLER_226_201 ();
 sky130_fd_sc_hs__fill_8 FILLER_226_204 ();
 sky130_fd_sc_hs__fill_1 FILLER_226_212 ();
 sky130_fd_sc_hs__fill_4 FILLER_226_255 ();
 sky130_fd_sc_hs__fill_2 FILLER_226_259 ();
 sky130_fd_sc_hs__fill_2 FILLER_226_262 ();
 sky130_fd_sc_hs__fill_1 FILLER_226_264 ();
 sky130_fd_sc_hs__fill_4 FILLER_226_270 ();
 sky130_fd_sc_hs__fill_1 FILLER_226_274 ();
 sky130_fd_sc_hs__fill_8 FILLER_226_288 ();
 sky130_fd_sc_hs__fill_8 FILLER_226_296 ();
 sky130_fd_sc_hs__fill_8 FILLER_226_304 ();
 sky130_fd_sc_hs__fill_4 FILLER_226_312 ();
 sky130_fd_sc_hs__fill_2 FILLER_226_316 ();
 sky130_fd_sc_hs__fill_1 FILLER_226_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_226_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_226_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_226_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_226_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_226_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_226_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_226_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_226_376 ();
 sky130_fd_sc_hs__fill_2 FILLER_226_378 ();
 sky130_fd_sc_hs__fill_1 FILLER_226_380 ();
 sky130_fd_sc_hs__fill_8 FILLER_226_383 ();
 sky130_fd_sc_hs__fill_8 FILLER_226_391 ();
 sky130_fd_sc_hs__fill_8 FILLER_226_399 ();
 sky130_fd_sc_hs__fill_8 FILLER_226_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_226_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_226_423 ();
 sky130_fd_sc_hs__fill_4 FILLER_226_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_226_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_226_444 ();
 sky130_fd_sc_hs__fill_4 FILLER_226_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_226_458 ();
 sky130_fd_sc_hs__fill_8 FILLER_226_466 ();
 sky130_fd_sc_hs__fill_8 FILLER_226_474 ();
 sky130_fd_sc_hs__fill_8 FILLER_226_482 ();
 sky130_fd_sc_hs__fill_2 FILLER_226_490 ();
 sky130_fd_sc_hs__fill_1 FILLER_226_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_226_494 ();
 sky130_fd_sc_hs__fill_4 FILLER_226_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_226_514 ();
 sky130_fd_sc_hs__fill_8 FILLER_226_522 ();
 sky130_fd_sc_hs__fill_8 FILLER_226_530 ();
 sky130_fd_sc_hs__fill_2 FILLER_226_538 ();
 sky130_fd_sc_hs__fill_8 FILLER_227_0 ();
 sky130_fd_sc_hs__fill_2 FILLER_227_8 ();
 sky130_fd_sc_hs__fill_1 FILLER_227_10 ();
 sky130_fd_sc_hs__fill_8 FILLER_227_19 ();
 sky130_fd_sc_hs__fill_8 FILLER_227_27 ();
 sky130_fd_sc_hs__fill_8 FILLER_227_35 ();
 sky130_fd_sc_hs__fill_2 FILLER_227_43 ();
 sky130_fd_sc_hs__fill_1 FILLER_227_57 ();
 sky130_fd_sc_hs__fill_8 FILLER_227_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_227_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_227_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_227_83 ();
 sky130_fd_sc_hs__fill_4 FILLER_227_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_227_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_227_125 ();
 sky130_fd_sc_hs__fill_8 FILLER_227_133 ();
 sky130_fd_sc_hs__fill_8 FILLER_227_141 ();
 sky130_fd_sc_hs__fill_2 FILLER_227_149 ();
 sky130_fd_sc_hs__fill_1 FILLER_227_151 ();
 sky130_fd_sc_hs__fill_1 FILLER_227_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_227_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_227_183 ();
 sky130_fd_sc_hs__fill_4 FILLER_227_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_227_208 ();
 sky130_fd_sc_hs__fill_8 FILLER_227_216 ();
 sky130_fd_sc_hs__fill_8 FILLER_227_224 ();
 sky130_fd_sc_hs__fill_4 FILLER_227_233 ();
 sky130_fd_sc_hs__fill_2 FILLER_227_237 ();
 sky130_fd_sc_hs__fill_8 FILLER_227_248 ();
 sky130_fd_sc_hs__fill_4 FILLER_227_256 ();
 sky130_fd_sc_hs__fill_1 FILLER_227_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_227_282 ();
 sky130_fd_sc_hs__fill_4 FILLER_227_291 ();
 sky130_fd_sc_hs__fill_4 FILLER_227_308 ();
 sky130_fd_sc_hs__fill_2 FILLER_227_312 ();
 sky130_fd_sc_hs__fill_1 FILLER_227_314 ();
 sky130_fd_sc_hs__fill_8 FILLER_227_335 ();
 sky130_fd_sc_hs__fill_4 FILLER_227_343 ();
 sky130_fd_sc_hs__fill_1 FILLER_227_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_227_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_227_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_227_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_227_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_227_383 ();
 sky130_fd_sc_hs__fill_8 FILLER_227_391 ();
 sky130_fd_sc_hs__fill_4 FILLER_227_399 ();
 sky130_fd_sc_hs__fill_2 FILLER_227_403 ();
 sky130_fd_sc_hs__fill_1 FILLER_227_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_227_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_227_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_227_423 ();
 sky130_fd_sc_hs__fill_8 FILLER_227_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_227_439 ();
 sky130_fd_sc_hs__fill_8 FILLER_227_447 ();
 sky130_fd_sc_hs__fill_1 FILLER_227_455 ();
 sky130_fd_sc_hs__fill_4 FILLER_227_458 ();
 sky130_fd_sc_hs__fill_2 FILLER_227_462 ();
 sky130_fd_sc_hs__fill_8 FILLER_227_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_227_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_227_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_227_489 ();
 sky130_fd_sc_hs__fill_1 FILLER_227_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_227_506 ();
 sky130_fd_sc_hs__fill_8 FILLER_227_514 ();
 sky130_fd_sc_hs__fill_8 FILLER_227_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_227_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_227_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_228_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_228_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_228_16 ();
 sky130_fd_sc_hs__fill_4 FILLER_228_24 ();
 sky130_fd_sc_hs__fill_1 FILLER_228_28 ();
 sky130_fd_sc_hs__fill_8 FILLER_228_30 ();
 sky130_fd_sc_hs__fill_4 FILLER_228_38 ();
 sky130_fd_sc_hs__fill_2 FILLER_228_42 ();
 sky130_fd_sc_hs__fill_8 FILLER_228_60 ();
 sky130_fd_sc_hs__fill_8 FILLER_228_68 ();
 sky130_fd_sc_hs__fill_8 FILLER_228_76 ();
 sky130_fd_sc_hs__fill_2 FILLER_228_84 ();
 sky130_fd_sc_hs__fill_1 FILLER_228_86 ();
 sky130_fd_sc_hs__fill_2 FILLER_228_88 ();
 sky130_fd_sc_hs__fill_1 FILLER_228_90 ();
 sky130_fd_sc_hs__fill_8 FILLER_228_133 ();
 sky130_fd_sc_hs__fill_4 FILLER_228_141 ();
 sky130_fd_sc_hs__fill_8 FILLER_228_146 ();
 sky130_fd_sc_hs__fill_2 FILLER_228_154 ();
 sky130_fd_sc_hs__fill_1 FILLER_228_156 ();
 sky130_fd_sc_hs__fill_4 FILLER_228_199 ();
 sky130_fd_sc_hs__fill_8 FILLER_228_204 ();
 sky130_fd_sc_hs__fill_8 FILLER_228_212 ();
 sky130_fd_sc_hs__fill_2 FILLER_228_220 ();
 sky130_fd_sc_hs__fill_8 FILLER_228_243 ();
 sky130_fd_sc_hs__fill_8 FILLER_228_251 ();
 sky130_fd_sc_hs__fill_2 FILLER_228_259 ();
 sky130_fd_sc_hs__fill_2 FILLER_228_280 ();
 sky130_fd_sc_hs__fill_1 FILLER_228_282 ();
 sky130_fd_sc_hs__fill_2 FILLER_228_304 ();
 sky130_fd_sc_hs__fill_1 FILLER_228_306 ();
 sky130_fd_sc_hs__fill_8 FILLER_228_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_228_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_228_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_228_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_228_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_228_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_228_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_228_376 ();
 sky130_fd_sc_hs__fill_2 FILLER_228_378 ();
 sky130_fd_sc_hs__fill_1 FILLER_228_380 ();
 sky130_fd_sc_hs__fill_8 FILLER_228_383 ();
 sky130_fd_sc_hs__fill_8 FILLER_228_391 ();
 sky130_fd_sc_hs__fill_8 FILLER_228_399 ();
 sky130_fd_sc_hs__fill_8 FILLER_228_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_228_415 ();
 sky130_fd_sc_hs__fill_8 FILLER_228_423 ();
 sky130_fd_sc_hs__fill_4 FILLER_228_431 ();
 sky130_fd_sc_hs__fill_8 FILLER_228_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_228_444 ();
 sky130_fd_sc_hs__fill_4 FILLER_228_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_228_458 ();
 sky130_fd_sc_hs__fill_8 FILLER_228_466 ();
 sky130_fd_sc_hs__fill_8 FILLER_228_474 ();
 sky130_fd_sc_hs__fill_8 FILLER_228_482 ();
 sky130_fd_sc_hs__fill_2 FILLER_228_490 ();
 sky130_fd_sc_hs__fill_1 FILLER_228_492 ();
 sky130_fd_sc_hs__fill_8 FILLER_228_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_228_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_228_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_228_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_228_526 ();
 sky130_fd_sc_hs__fill_4 FILLER_228_534 ();
 sky130_fd_sc_hs__fill_2 FILLER_228_538 ();
 sky130_fd_sc_hs__fill_8 FILLER_229_0 ();
 sky130_fd_sc_hs__fill_4 FILLER_229_8 ();
 sky130_fd_sc_hs__fill_1 FILLER_229_12 ();
 sky130_fd_sc_hs__fill_8 FILLER_229_21 ();
 sky130_fd_sc_hs__fill_8 FILLER_229_29 ();
 sky130_fd_sc_hs__fill_8 FILLER_229_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_229_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_229_117 ();
 sky130_fd_sc_hs__fill_4 FILLER_229_125 ();
 sky130_fd_sc_hs__fill_2 FILLER_229_129 ();
 sky130_fd_sc_hs__fill_1 FILLER_229_173 ();
 sky130_fd_sc_hs__fill_8 FILLER_229_196 ();
 sky130_fd_sc_hs__fill_4 FILLER_229_204 ();
 sky130_fd_sc_hs__fill_1 FILLER_229_208 ();
 sky130_fd_sc_hs__fill_8 FILLER_229_221 ();
 sky130_fd_sc_hs__fill_2 FILLER_229_229 ();
 sky130_fd_sc_hs__fill_1 FILLER_229_231 ();
 sky130_fd_sc_hs__fill_4 FILLER_229_233 ();
 sky130_fd_sc_hs__fill_2 FILLER_229_237 ();
 sky130_fd_sc_hs__fill_1 FILLER_229_239 ();
 sky130_fd_sc_hs__fill_1 FILLER_229_289 ();
 sky130_fd_sc_hs__fill_2 FILLER_229_291 ();
 sky130_fd_sc_hs__fill_1 FILLER_229_293 ();
 sky130_fd_sc_hs__fill_8 FILLER_229_326 ();
 sky130_fd_sc_hs__fill_8 FILLER_229_334 ();
 sky130_fd_sc_hs__fill_4 FILLER_229_342 ();
 sky130_fd_sc_hs__fill_2 FILLER_229_346 ();
 sky130_fd_sc_hs__fill_8 FILLER_229_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_229_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_229_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_229_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_229_383 ();
 sky130_fd_sc_hs__fill_8 FILLER_229_391 ();
 sky130_fd_sc_hs__fill_4 FILLER_229_399 ();
 sky130_fd_sc_hs__fill_2 FILLER_229_403 ();
 sky130_fd_sc_hs__fill_1 FILLER_229_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_229_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_229_417 ();
 sky130_fd_sc_hs__fill_8 FILLER_229_425 ();
 sky130_fd_sc_hs__fill_8 FILLER_229_433 ();
 sky130_fd_sc_hs__fill_8 FILLER_229_441 ();
 sky130_fd_sc_hs__fill_4 FILLER_229_449 ();
 sky130_fd_sc_hs__fill_1 FILLER_229_455 ();
 sky130_fd_sc_hs__fill_4 FILLER_229_458 ();
 sky130_fd_sc_hs__fill_2 FILLER_229_462 ();
 sky130_fd_sc_hs__fill_8 FILLER_229_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_229_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_229_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_229_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_229_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_229_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_229_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_229_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_229_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_229_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_229_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_230_0 ();
 sky130_fd_sc_hs__fill_1 FILLER_230_8 ();
 sky130_fd_sc_hs__fill_4 FILLER_230_25 ();
 sky130_fd_sc_hs__fill_8 FILLER_230_30 ();
 sky130_fd_sc_hs__fill_8 FILLER_230_38 ();
 sky130_fd_sc_hs__fill_1 FILLER_230_46 ();
 sky130_fd_sc_hs__fill_8 FILLER_230_68 ();
 sky130_fd_sc_hs__fill_8 FILLER_230_76 ();
 sky130_fd_sc_hs__fill_2 FILLER_230_84 ();
 sky130_fd_sc_hs__fill_1 FILLER_230_86 ();
 sky130_fd_sc_hs__fill_8 FILLER_230_129 ();
 sky130_fd_sc_hs__fill_8 FILLER_230_137 ();
 sky130_fd_sc_hs__fill_8 FILLER_230_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_230_154 ();
 sky130_fd_sc_hs__fill_8 FILLER_230_162 ();
 sky130_fd_sc_hs__fill_8 FILLER_230_170 ();
 sky130_fd_sc_hs__fill_4 FILLER_230_178 ();
 sky130_fd_sc_hs__fill_1 FILLER_230_182 ();
 sky130_fd_sc_hs__fill_8 FILLER_230_204 ();
 sky130_fd_sc_hs__fill_4 FILLER_230_212 ();
 sky130_fd_sc_hs__fill_2 FILLER_230_216 ();
 sky130_fd_sc_hs__fill_1 FILLER_230_218 ();
 sky130_fd_sc_hs__fill_8 FILLER_230_248 ();
 sky130_fd_sc_hs__fill_4 FILLER_230_256 ();
 sky130_fd_sc_hs__fill_1 FILLER_230_260 ();
 sky130_fd_sc_hs__fill_8 FILLER_230_271 ();
 sky130_fd_sc_hs__fill_8 FILLER_230_292 ();
 sky130_fd_sc_hs__fill_8 FILLER_230_300 ();
 sky130_fd_sc_hs__fill_8 FILLER_230_308 ();
 sky130_fd_sc_hs__fill_2 FILLER_230_316 ();
 sky130_fd_sc_hs__fill_1 FILLER_230_318 ();
 sky130_fd_sc_hs__fill_8 FILLER_230_320 ();
 sky130_fd_sc_hs__fill_8 FILLER_230_328 ();
 sky130_fd_sc_hs__fill_8 FILLER_230_336 ();
 sky130_fd_sc_hs__fill_8 FILLER_230_344 ();
 sky130_fd_sc_hs__fill_8 FILLER_230_352 ();
 sky130_fd_sc_hs__fill_8 FILLER_230_360 ();
 sky130_fd_sc_hs__fill_8 FILLER_230_368 ();
 sky130_fd_sc_hs__fill_1 FILLER_230_376 ();
 sky130_fd_sc_hs__fill_2 FILLER_230_378 ();
 sky130_fd_sc_hs__fill_1 FILLER_230_380 ();
 sky130_fd_sc_hs__fill_8 FILLER_230_383 ();
 sky130_fd_sc_hs__fill_8 FILLER_230_391 ();
 sky130_fd_sc_hs__fill_8 FILLER_230_399 ();
 sky130_fd_sc_hs__fill_8 FILLER_230_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_230_417 ();
 sky130_fd_sc_hs__fill_8 FILLER_230_425 ();
 sky130_fd_sc_hs__fill_2 FILLER_230_433 ();
 sky130_fd_sc_hs__fill_8 FILLER_230_436 ();
 sky130_fd_sc_hs__fill_8 FILLER_230_444 ();
 sky130_fd_sc_hs__fill_1 FILLER_230_452 ();
 sky130_fd_sc_hs__fill_8 FILLER_230_461 ();
 sky130_fd_sc_hs__fill_8 FILLER_230_469 ();
 sky130_fd_sc_hs__fill_8 FILLER_230_477 ();
 sky130_fd_sc_hs__fill_8 FILLER_230_485 ();
 sky130_fd_sc_hs__fill_8 FILLER_230_494 ();
 sky130_fd_sc_hs__fill_8 FILLER_230_502 ();
 sky130_fd_sc_hs__fill_8 FILLER_230_510 ();
 sky130_fd_sc_hs__fill_8 FILLER_230_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_230_526 ();
 sky130_fd_sc_hs__fill_4 FILLER_230_534 ();
 sky130_fd_sc_hs__fill_2 FILLER_230_538 ();
 sky130_fd_sc_hs__fill_8 FILLER_231_0 ();
 sky130_fd_sc_hs__fill_8 FILLER_231_8 ();
 sky130_fd_sc_hs__fill_8 FILLER_231_16 ();
 sky130_fd_sc_hs__fill_8 FILLER_231_24 ();
 sky130_fd_sc_hs__fill_4 FILLER_231_32 ();
 sky130_fd_sc_hs__fill_1 FILLER_231_36 ();
 sky130_fd_sc_hs__fill_4 FILLER_231_45 ();
 sky130_fd_sc_hs__fill_1 FILLER_231_49 ();
 sky130_fd_sc_hs__fill_8 FILLER_231_59 ();
 sky130_fd_sc_hs__fill_8 FILLER_231_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_231_75 ();
 sky130_fd_sc_hs__fill_8 FILLER_231_83 ();
 sky130_fd_sc_hs__fill_8 FILLER_231_91 ();
 sky130_fd_sc_hs__fill_8 FILLER_231_99 ();
 sky130_fd_sc_hs__fill_8 FILLER_231_107 ();
 sky130_fd_sc_hs__fill_1 FILLER_231_115 ();
 sky130_fd_sc_hs__fill_1 FILLER_231_117 ();
 sky130_fd_sc_hs__fill_2 FILLER_231_126 ();
 sky130_fd_sc_hs__fill_1 FILLER_231_128 ();
 sky130_fd_sc_hs__fill_8 FILLER_231_137 ();
 sky130_fd_sc_hs__fill_1 FILLER_231_145 ();
 sky130_fd_sc_hs__fill_8 FILLER_231_162 ();
 sky130_fd_sc_hs__fill_4 FILLER_231_170 ();
 sky130_fd_sc_hs__fill_8 FILLER_231_175 ();
 sky130_fd_sc_hs__fill_8 FILLER_231_183 ();
 sky130_fd_sc_hs__fill_8 FILLER_231_191 ();
 sky130_fd_sc_hs__fill_8 FILLER_231_199 ();
 sky130_fd_sc_hs__fill_2 FILLER_231_207 ();
 sky130_fd_sc_hs__fill_8 FILLER_231_217 ();
 sky130_fd_sc_hs__fill_4 FILLER_231_225 ();
 sky130_fd_sc_hs__fill_2 FILLER_231_229 ();
 sky130_fd_sc_hs__fill_1 FILLER_231_231 ();
 sky130_fd_sc_hs__fill_8 FILLER_231_233 ();
 sky130_fd_sc_hs__fill_8 FILLER_231_241 ();
 sky130_fd_sc_hs__fill_8 FILLER_231_249 ();
 sky130_fd_sc_hs__fill_8 FILLER_231_257 ();
 sky130_fd_sc_hs__fill_8 FILLER_231_265 ();
 sky130_fd_sc_hs__fill_8 FILLER_231_273 ();
 sky130_fd_sc_hs__fill_1 FILLER_231_281 ();
 sky130_fd_sc_hs__fill_2 FILLER_231_291 ();
 sky130_fd_sc_hs__fill_8 FILLER_231_301 ();
 sky130_fd_sc_hs__fill_8 FILLER_231_309 ();
 sky130_fd_sc_hs__fill_8 FILLER_231_317 ();
 sky130_fd_sc_hs__fill_4 FILLER_231_325 ();
 sky130_fd_sc_hs__fill_8 FILLER_231_337 ();
 sky130_fd_sc_hs__fill_2 FILLER_231_345 ();
 sky130_fd_sc_hs__fill_1 FILLER_231_347 ();
 sky130_fd_sc_hs__fill_8 FILLER_231_349 ();
 sky130_fd_sc_hs__fill_8 FILLER_231_357 ();
 sky130_fd_sc_hs__fill_8 FILLER_231_365 ();
 sky130_fd_sc_hs__fill_8 FILLER_231_373 ();
 sky130_fd_sc_hs__fill_8 FILLER_231_383 ();
 sky130_fd_sc_hs__fill_8 FILLER_231_391 ();
 sky130_fd_sc_hs__fill_4 FILLER_231_399 ();
 sky130_fd_sc_hs__fill_2 FILLER_231_403 ();
 sky130_fd_sc_hs__fill_1 FILLER_231_405 ();
 sky130_fd_sc_hs__fill_8 FILLER_231_407 ();
 sky130_fd_sc_hs__fill_8 FILLER_231_425 ();
 sky130_fd_sc_hs__fill_8 FILLER_231_433 ();
 sky130_fd_sc_hs__fill_8 FILLER_231_441 ();
 sky130_fd_sc_hs__fill_4 FILLER_231_449 ();
 sky130_fd_sc_hs__fill_1 FILLER_231_455 ();
 sky130_fd_sc_hs__fill_4 FILLER_231_458 ();
 sky130_fd_sc_hs__fill_2 FILLER_231_462 ();
 sky130_fd_sc_hs__fill_8 FILLER_231_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_231_473 ();
 sky130_fd_sc_hs__fill_8 FILLER_231_481 ();
 sky130_fd_sc_hs__fill_8 FILLER_231_489 ();
 sky130_fd_sc_hs__fill_8 FILLER_231_497 ();
 sky130_fd_sc_hs__fill_8 FILLER_231_505 ();
 sky130_fd_sc_hs__fill_8 FILLER_231_513 ();
 sky130_fd_sc_hs__fill_1 FILLER_231_521 ();
 sky130_fd_sc_hs__fill_8 FILLER_231_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_231_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_231_539 ();
 sky130_fd_sc_hs__fill_8 FILLER_232_0 ();
 sky130_fd_sc_hs__fill_4 FILLER_232_8 ();
 sky130_fd_sc_hs__fill_1 FILLER_232_12 ();
 sky130_fd_sc_hs__fill_8 FILLER_232_21 ();
 sky130_fd_sc_hs__fill_2 FILLER_232_30 ();
 sky130_fd_sc_hs__fill_2 FILLER_232_48 ();
 sky130_fd_sc_hs__fill_4 FILLER_232_67 ();
 sky130_fd_sc_hs__fill_8 FILLER_232_79 ();
 sky130_fd_sc_hs__fill_2 FILLER_232_88 ();
 sky130_fd_sc_hs__fill_8 FILLER_232_98 ();
 sky130_fd_sc_hs__fill_8 FILLER_232_106 ();
 sky130_fd_sc_hs__fill_2 FILLER_232_114 ();
 sky130_fd_sc_hs__fill_2 FILLER_232_117 ();
 sky130_fd_sc_hs__fill_8 FILLER_232_127 ();
 sky130_fd_sc_hs__fill_2 FILLER_232_135 ();
 sky130_fd_sc_hs__fill_4 FILLER_232_146 ();
 sky130_fd_sc_hs__fill_8 FILLER_232_175 ();
 sky130_fd_sc_hs__fill_4 FILLER_232_183 ();
 sky130_fd_sc_hs__fill_1 FILLER_232_204 ();
 sky130_fd_sc_hs__fill_1 FILLER_232_213 ();
 sky130_fd_sc_hs__fill_8 FILLER_232_222 ();
 sky130_fd_sc_hs__fill_2 FILLER_232_230 ();
 sky130_fd_sc_hs__fill_1 FILLER_232_241 ();
 sky130_fd_sc_hs__fill_1 FILLER_232_250 ();
 sky130_fd_sc_hs__fill_2 FILLER_232_259 ();
 sky130_fd_sc_hs__fill_8 FILLER_232_262 ();
 sky130_fd_sc_hs__fill_4 FILLER_232_270 ();
 sky130_fd_sc_hs__fill_4 FILLER_232_299 ();
 sky130_fd_sc_hs__fill_1 FILLER_232_320 ();
 sky130_fd_sc_hs__fill_2 FILLER_232_337 ();
 sky130_fd_sc_hs__fill_1 FILLER_232_339 ();
 sky130_fd_sc_hs__fill_4 FILLER_232_365 ();
 sky130_fd_sc_hs__fill_2 FILLER_232_378 ();
 sky130_fd_sc_hs__fill_1 FILLER_232_380 ();
 sky130_fd_sc_hs__fill_1 FILLER_232_389 ();
 sky130_fd_sc_hs__fill_4 FILLER_232_431 ();
 sky130_fd_sc_hs__fill_4 FILLER_232_436 ();
 sky130_fd_sc_hs__fill_4 FILLER_232_465 ();
 sky130_fd_sc_hs__fill_8 FILLER_232_477 ();
 sky130_fd_sc_hs__fill_4 FILLER_232_518 ();
 sky130_fd_sc_hs__fill_8 FILLER_232_523 ();
 sky130_fd_sc_hs__fill_8 FILLER_232_531 ();
 sky130_fd_sc_hs__fill_1 FILLER_232_539 ();
endmodule
