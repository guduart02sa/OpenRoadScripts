VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 1000 ;
END UNITS

VIA ibex_wb_stage_via2_3_1600_480_1_5_320_320
  VIARULE M1M2_PR ;
  CUTSIZE 0.15 0.15 ;
  LAYERS met1 via met2 ;
  CUTSPACING 0.17 0.17 ;
  ENCLOSURE 0.085 0.165 0.055 0.085 ;
  ROWCOL 1 5 ;
END ibex_wb_stage_via2_3_1600_480_1_5_320_320

VIA ibex_wb_stage_via3_4_1600_480_1_4_400_400
  VIARULE M2M3_PR ;
  CUTSIZE 0.2 0.2 ;
  LAYERS met2 via2 met3 ;
  CUTSPACING 0.2 0.2 ;
  ENCLOSURE 0.04 0.085 0.065 0.065 ;
  ROWCOL 1 4 ;
END ibex_wb_stage_via3_4_1600_480_1_4_400_400

VIA ibex_wb_stage_via4_5_1600_480_1_4_400_400
  VIARULE M3M4_PR ;
  CUTSIZE 0.2 0.2 ;
  LAYERS met3 via3 met4 ;
  CUTSPACING 0.2 0.2 ;
  ENCLOSURE 0.09 0.06 0.1 0.065 ;
  ROWCOL 1 4 ;
END ibex_wb_stage_via4_5_1600_480_1_4_400_400

VIA ibex_wb_stage_via5_6_1600_1600_1_1_1600_1600
  VIARULE M4M5_PR ;
  CUTSIZE 0.8 0.8 ;
  LAYERS met4 via4 met5 ;
  CUTSPACING 0.8 0.8 ;
  ENCLOSURE 0.4 0.19 0.31 0.4 ;
END ibex_wb_stage_via5_6_1600_1600_1_1_1600_1600

MACRO ibex_wb_stage
  FOREIGN ibex_wb_stage 0 0 ;
  CLASS BLOCK ;
  SIZE 58.02 BY 170.065 ;
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      LAYER met5 ;
        RECT  27.72 165.12 56.46 166.72 ;
        RECT  27.72 137.92 56.46 139.52 ;
        RECT  27.72 110.72 56.46 112.32 ;
        RECT  27.72 83.52 56.46 85.12 ;
        RECT  27.72 56.32 56.46 57.92 ;
        RECT  27.72 29.12 56.46 30.72 ;
      LAYER met4 ;
        RECT  54.86 5.2 56.46 168.88 ;
        RECT  27.72 5.2 29.32 168.88 ;
      LAYER met1 ;
        RECT  1.38 168.4 56.58 168.88 ;
        RECT  1.38 162.96 56.58 163.44 ;
        RECT  1.38 157.52 56.58 158 ;
        RECT  1.38 152.08 56.58 152.56 ;
        RECT  1.38 146.64 56.58 147.12 ;
        RECT  1.38 141.2 56.58 141.68 ;
        RECT  1.38 135.76 56.58 136.24 ;
        RECT  1.38 130.32 56.58 130.8 ;
        RECT  1.38 124.88 56.58 125.36 ;
        RECT  1.38 119.44 56.58 119.92 ;
        RECT  1.38 114 56.58 114.48 ;
        RECT  1.38 108.56 56.58 109.04 ;
        RECT  1.38 103.12 56.58 103.6 ;
        RECT  1.38 97.68 56.58 98.16 ;
        RECT  1.38 92.24 56.58 92.72 ;
        RECT  1.38 86.8 56.58 87.28 ;
        RECT  1.38 81.36 56.58 81.84 ;
        RECT  1.38 75.92 56.58 76.4 ;
        RECT  1.38 70.48 56.58 70.96 ;
        RECT  1.38 65.04 56.58 65.52 ;
        RECT  1.38 59.6 56.58 60.08 ;
        RECT  1.38 54.16 56.58 54.64 ;
        RECT  1.38 48.72 56.58 49.2 ;
        RECT  1.38 43.28 56.58 43.76 ;
        RECT  1.38 37.84 56.58 38.32 ;
        RECT  1.38 32.4 56.58 32.88 ;
        RECT  1.38 26.96 56.58 27.44 ;
        RECT  1.38 21.52 56.58 22 ;
        RECT  1.38 16.08 56.58 16.56 ;
        RECT  1.38 10.64 56.58 11.12 ;
        RECT  1.38 5.2 56.58 5.68 ;
      VIA 55.66 165.92 ibex_wb_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 138.72 ibex_wb_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 111.52 ibex_wb_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 84.32 ibex_wb_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 57.12 ibex_wb_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 29.92 ibex_wb_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 165.92 ibex_wb_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 138.72 ibex_wb_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 111.52 ibex_wb_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 84.32 ibex_wb_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 57.12 ibex_wb_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 29.92 ibex_wb_stage_via5_6_1600_1600_1_1_1600_1600 ;
      LAYER met3 ;
        RECT  54.87 168.475 56.45 168.805 ;
      VIA 55.66 168.64 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 168.455 56.43 168.825 ;
      VIA 55.66 168.64 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 168.64 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 163.035 56.45 163.365 ;
      VIA 55.66 163.2 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 163.015 56.43 163.385 ;
      VIA 55.66 163.2 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 163.2 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 157.595 56.45 157.925 ;
      VIA 55.66 157.76 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 157.575 56.43 157.945 ;
      VIA 55.66 157.76 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 157.76 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 152.155 56.45 152.485 ;
      VIA 55.66 152.32 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 152.135 56.43 152.505 ;
      VIA 55.66 152.32 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 152.32 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 146.715 56.45 147.045 ;
      VIA 55.66 146.88 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 146.695 56.43 147.065 ;
      VIA 55.66 146.88 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 146.88 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 141.275 56.45 141.605 ;
      VIA 55.66 141.44 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 141.255 56.43 141.625 ;
      VIA 55.66 141.44 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 141.44 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 135.835 56.45 136.165 ;
      VIA 55.66 136 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 135.815 56.43 136.185 ;
      VIA 55.66 136 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 136 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 130.395 56.45 130.725 ;
      VIA 55.66 130.56 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 130.375 56.43 130.745 ;
      VIA 55.66 130.56 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 130.56 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 124.955 56.45 125.285 ;
      VIA 55.66 125.12 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 124.935 56.43 125.305 ;
      VIA 55.66 125.12 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 125.12 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 119.515 56.45 119.845 ;
      VIA 55.66 119.68 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 119.495 56.43 119.865 ;
      VIA 55.66 119.68 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 119.68 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 114.075 56.45 114.405 ;
      VIA 55.66 114.24 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 114.055 56.43 114.425 ;
      VIA 55.66 114.24 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 114.24 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 108.635 56.45 108.965 ;
      VIA 55.66 108.8 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 108.615 56.43 108.985 ;
      VIA 55.66 108.8 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 108.8 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 103.195 56.45 103.525 ;
      VIA 55.66 103.36 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 103.175 56.43 103.545 ;
      VIA 55.66 103.36 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 103.36 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 97.755 56.45 98.085 ;
      VIA 55.66 97.92 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 97.735 56.43 98.105 ;
      VIA 55.66 97.92 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 97.92 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 92.315 56.45 92.645 ;
      VIA 55.66 92.48 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 92.295 56.43 92.665 ;
      VIA 55.66 92.48 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 92.48 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 86.875 56.45 87.205 ;
      VIA 55.66 87.04 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 86.855 56.43 87.225 ;
      VIA 55.66 87.04 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 87.04 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 81.435 56.45 81.765 ;
      VIA 55.66 81.6 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 81.415 56.43 81.785 ;
      VIA 55.66 81.6 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 81.6 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 75.995 56.45 76.325 ;
      VIA 55.66 76.16 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 75.975 56.43 76.345 ;
      VIA 55.66 76.16 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 76.16 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 70.555 56.45 70.885 ;
      VIA 55.66 70.72 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 70.535 56.43 70.905 ;
      VIA 55.66 70.72 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 70.72 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 65.115 56.45 65.445 ;
      VIA 55.66 65.28 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 65.095 56.43 65.465 ;
      VIA 55.66 65.28 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 65.28 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 59.675 56.45 60.005 ;
      VIA 55.66 59.84 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 59.655 56.43 60.025 ;
      VIA 55.66 59.84 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 59.84 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 54.235 56.45 54.565 ;
      VIA 55.66 54.4 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 54.215 56.43 54.585 ;
      VIA 55.66 54.4 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 54.4 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 48.795 56.45 49.125 ;
      VIA 55.66 48.96 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 48.775 56.43 49.145 ;
      VIA 55.66 48.96 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 48.96 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 43.355 56.45 43.685 ;
      VIA 55.66 43.52 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 43.335 56.43 43.705 ;
      VIA 55.66 43.52 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 43.52 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 37.915 56.45 38.245 ;
      VIA 55.66 38.08 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 37.895 56.43 38.265 ;
      VIA 55.66 38.08 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 38.08 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 32.475 56.45 32.805 ;
      VIA 55.66 32.64 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 32.455 56.43 32.825 ;
      VIA 55.66 32.64 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 32.64 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 27.035 56.45 27.365 ;
      VIA 55.66 27.2 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 27.015 56.43 27.385 ;
      VIA 55.66 27.2 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 27.2 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 21.595 56.45 21.925 ;
      VIA 55.66 21.76 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 21.575 56.43 21.945 ;
      VIA 55.66 21.76 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 21.76 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 16.155 56.45 16.485 ;
      VIA 55.66 16.32 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 16.135 56.43 16.505 ;
      VIA 55.66 16.32 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 16.32 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 10.715 56.45 11.045 ;
      VIA 55.66 10.88 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 10.695 56.43 11.065 ;
      VIA 55.66 10.88 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 10.88 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 5.275 56.45 5.605 ;
      VIA 55.66 5.44 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 5.255 56.43 5.625 ;
      VIA 55.66 5.44 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 5.44 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 168.475 29.31 168.805 ;
      VIA 28.52 168.64 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 168.455 29.29 168.825 ;
      VIA 28.52 168.64 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 168.64 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 163.035 29.31 163.365 ;
      VIA 28.52 163.2 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 163.015 29.29 163.385 ;
      VIA 28.52 163.2 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 163.2 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 157.595 29.31 157.925 ;
      VIA 28.52 157.76 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 157.575 29.29 157.945 ;
      VIA 28.52 157.76 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 157.76 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 152.155 29.31 152.485 ;
      VIA 28.52 152.32 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 152.135 29.29 152.505 ;
      VIA 28.52 152.32 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 152.32 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 146.715 29.31 147.045 ;
      VIA 28.52 146.88 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 146.695 29.29 147.065 ;
      VIA 28.52 146.88 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 146.88 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 141.275 29.31 141.605 ;
      VIA 28.52 141.44 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 141.255 29.29 141.625 ;
      VIA 28.52 141.44 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 141.44 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 135.835 29.31 136.165 ;
      VIA 28.52 136 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 135.815 29.29 136.185 ;
      VIA 28.52 136 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 136 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 130.395 29.31 130.725 ;
      VIA 28.52 130.56 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 130.375 29.29 130.745 ;
      VIA 28.52 130.56 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 130.56 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 124.955 29.31 125.285 ;
      VIA 28.52 125.12 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 124.935 29.29 125.305 ;
      VIA 28.52 125.12 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 125.12 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 119.515 29.31 119.845 ;
      VIA 28.52 119.68 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 119.495 29.29 119.865 ;
      VIA 28.52 119.68 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 119.68 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 114.075 29.31 114.405 ;
      VIA 28.52 114.24 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 114.055 29.29 114.425 ;
      VIA 28.52 114.24 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 114.24 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 108.635 29.31 108.965 ;
      VIA 28.52 108.8 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 108.615 29.29 108.985 ;
      VIA 28.52 108.8 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 108.8 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 103.195 29.31 103.525 ;
      VIA 28.52 103.36 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 103.175 29.29 103.545 ;
      VIA 28.52 103.36 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 103.36 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 97.755 29.31 98.085 ;
      VIA 28.52 97.92 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 97.735 29.29 98.105 ;
      VIA 28.52 97.92 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 97.92 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 92.315 29.31 92.645 ;
      VIA 28.52 92.48 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 92.295 29.29 92.665 ;
      VIA 28.52 92.48 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 92.48 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 86.875 29.31 87.205 ;
      VIA 28.52 87.04 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 86.855 29.29 87.225 ;
      VIA 28.52 87.04 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 87.04 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 81.435 29.31 81.765 ;
      VIA 28.52 81.6 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 81.415 29.29 81.785 ;
      VIA 28.52 81.6 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 81.6 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 75.995 29.31 76.325 ;
      VIA 28.52 76.16 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 75.975 29.29 76.345 ;
      VIA 28.52 76.16 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 76.16 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 70.555 29.31 70.885 ;
      VIA 28.52 70.72 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 70.535 29.29 70.905 ;
      VIA 28.52 70.72 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 70.72 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 65.115 29.31 65.445 ;
      VIA 28.52 65.28 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 65.095 29.29 65.465 ;
      VIA 28.52 65.28 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 65.28 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 59.675 29.31 60.005 ;
      VIA 28.52 59.84 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 59.655 29.29 60.025 ;
      VIA 28.52 59.84 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 59.84 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 54.235 29.31 54.565 ;
      VIA 28.52 54.4 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 54.215 29.29 54.585 ;
      VIA 28.52 54.4 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 54.4 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 48.795 29.31 49.125 ;
      VIA 28.52 48.96 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 48.775 29.29 49.145 ;
      VIA 28.52 48.96 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 48.96 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 43.355 29.31 43.685 ;
      VIA 28.52 43.52 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 43.335 29.29 43.705 ;
      VIA 28.52 43.52 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 43.52 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 37.915 29.31 38.245 ;
      VIA 28.52 38.08 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 37.895 29.29 38.265 ;
      VIA 28.52 38.08 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 38.08 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 32.475 29.31 32.805 ;
      VIA 28.52 32.64 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 32.455 29.29 32.825 ;
      VIA 28.52 32.64 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 32.64 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 27.035 29.31 27.365 ;
      VIA 28.52 27.2 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 27.015 29.29 27.385 ;
      VIA 28.52 27.2 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 27.2 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 21.595 29.31 21.925 ;
      VIA 28.52 21.76 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 21.575 29.29 21.945 ;
      VIA 28.52 21.76 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 21.76 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 16.155 29.31 16.485 ;
      VIA 28.52 16.32 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 16.135 29.29 16.505 ;
      VIA 28.52 16.32 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 16.32 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 10.715 29.31 11.045 ;
      VIA 28.52 10.88 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 10.695 29.29 11.065 ;
      VIA 28.52 10.88 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 10.88 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 5.275 29.31 5.605 ;
      VIA 28.52 5.44 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 5.255 29.29 5.625 ;
      VIA 28.52 5.44 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 5.44 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      LAYER met5 ;
        RECT  14.15 151.52 42.89 153.12 ;
        RECT  14.15 124.32 42.89 125.92 ;
        RECT  14.15 97.12 42.89 98.72 ;
        RECT  14.15 69.92 42.89 71.52 ;
        RECT  14.15 42.72 42.89 44.32 ;
        RECT  14.15 15.52 42.89 17.12 ;
      LAYER met4 ;
        RECT  41.29 2.48 42.89 166.16 ;
        RECT  14.15 2.48 15.75 166.16 ;
      LAYER met1 ;
        RECT  1.38 165.68 56.58 166.16 ;
        RECT  1.38 160.24 56.58 160.72 ;
        RECT  1.38 154.8 56.58 155.28 ;
        RECT  1.38 149.36 56.58 149.84 ;
        RECT  1.38 143.92 56.58 144.4 ;
        RECT  1.38 138.48 56.58 138.96 ;
        RECT  1.38 133.04 56.58 133.52 ;
        RECT  1.38 127.6 56.58 128.08 ;
        RECT  1.38 122.16 56.58 122.64 ;
        RECT  1.38 116.72 56.58 117.2 ;
        RECT  1.38 111.28 56.58 111.76 ;
        RECT  1.38 105.84 56.58 106.32 ;
        RECT  1.38 100.4 56.58 100.88 ;
        RECT  1.38 94.96 56.58 95.44 ;
        RECT  1.38 89.52 56.58 90 ;
        RECT  1.38 84.08 56.58 84.56 ;
        RECT  1.38 78.64 56.58 79.12 ;
        RECT  1.38 73.2 56.58 73.68 ;
        RECT  1.38 67.76 56.58 68.24 ;
        RECT  1.38 62.32 56.58 62.8 ;
        RECT  1.38 56.88 56.58 57.36 ;
        RECT  1.38 51.44 56.58 51.92 ;
        RECT  1.38 46 56.58 46.48 ;
        RECT  1.38 40.56 56.58 41.04 ;
        RECT  1.38 35.12 56.58 35.6 ;
        RECT  1.38 29.68 56.58 30.16 ;
        RECT  1.38 24.24 56.58 24.72 ;
        RECT  1.38 18.8 56.58 19.28 ;
        RECT  1.38 13.36 56.58 13.84 ;
        RECT  1.38 7.92 56.58 8.4 ;
        RECT  1.38 2.48 56.58 2.96 ;
      VIA 42.09 152.32 ibex_wb_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 125.12 ibex_wb_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 97.92 ibex_wb_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 70.72 ibex_wb_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 43.52 ibex_wb_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 16.32 ibex_wb_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 152.32 ibex_wb_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 125.12 ibex_wb_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 97.92 ibex_wb_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 70.72 ibex_wb_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 43.52 ibex_wb_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 16.32 ibex_wb_stage_via5_6_1600_1600_1_1_1600_1600 ;
      LAYER met3 ;
        RECT  41.3 165.755 42.88 166.085 ;
      VIA 42.09 165.92 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 165.735 42.86 166.105 ;
      VIA 42.09 165.92 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 165.92 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 160.315 42.88 160.645 ;
      VIA 42.09 160.48 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 160.295 42.86 160.665 ;
      VIA 42.09 160.48 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 160.48 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 154.875 42.88 155.205 ;
      VIA 42.09 155.04 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 154.855 42.86 155.225 ;
      VIA 42.09 155.04 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 155.04 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 149.435 42.88 149.765 ;
      VIA 42.09 149.6 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 149.415 42.86 149.785 ;
      VIA 42.09 149.6 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 149.6 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 143.995 42.88 144.325 ;
      VIA 42.09 144.16 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 143.975 42.86 144.345 ;
      VIA 42.09 144.16 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 144.16 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 138.555 42.88 138.885 ;
      VIA 42.09 138.72 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 138.535 42.86 138.905 ;
      VIA 42.09 138.72 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 138.72 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 133.115 42.88 133.445 ;
      VIA 42.09 133.28 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 133.095 42.86 133.465 ;
      VIA 42.09 133.28 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 133.28 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 127.675 42.88 128.005 ;
      VIA 42.09 127.84 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 127.655 42.86 128.025 ;
      VIA 42.09 127.84 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 127.84 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 122.235 42.88 122.565 ;
      VIA 42.09 122.4 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 122.215 42.86 122.585 ;
      VIA 42.09 122.4 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 122.4 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 116.795 42.88 117.125 ;
      VIA 42.09 116.96 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 116.775 42.86 117.145 ;
      VIA 42.09 116.96 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 116.96 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 111.355 42.88 111.685 ;
      VIA 42.09 111.52 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 111.335 42.86 111.705 ;
      VIA 42.09 111.52 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 111.52 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 105.915 42.88 106.245 ;
      VIA 42.09 106.08 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 105.895 42.86 106.265 ;
      VIA 42.09 106.08 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 106.08 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 100.475 42.88 100.805 ;
      VIA 42.09 100.64 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 100.455 42.86 100.825 ;
      VIA 42.09 100.64 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 100.64 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 95.035 42.88 95.365 ;
      VIA 42.09 95.2 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 95.015 42.86 95.385 ;
      VIA 42.09 95.2 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 95.2 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 89.595 42.88 89.925 ;
      VIA 42.09 89.76 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 89.575 42.86 89.945 ;
      VIA 42.09 89.76 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 89.76 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 84.155 42.88 84.485 ;
      VIA 42.09 84.32 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 84.135 42.86 84.505 ;
      VIA 42.09 84.32 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 84.32 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 78.715 42.88 79.045 ;
      VIA 42.09 78.88 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 78.695 42.86 79.065 ;
      VIA 42.09 78.88 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 78.88 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 73.275 42.88 73.605 ;
      VIA 42.09 73.44 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 73.255 42.86 73.625 ;
      VIA 42.09 73.44 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 73.44 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 67.835 42.88 68.165 ;
      VIA 42.09 68 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 67.815 42.86 68.185 ;
      VIA 42.09 68 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 68 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 62.395 42.88 62.725 ;
      VIA 42.09 62.56 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 62.375 42.86 62.745 ;
      VIA 42.09 62.56 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 62.56 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 56.955 42.88 57.285 ;
      VIA 42.09 57.12 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 56.935 42.86 57.305 ;
      VIA 42.09 57.12 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 57.12 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 51.515 42.88 51.845 ;
      VIA 42.09 51.68 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 51.495 42.86 51.865 ;
      VIA 42.09 51.68 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 51.68 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 46.075 42.88 46.405 ;
      VIA 42.09 46.24 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 46.055 42.86 46.425 ;
      VIA 42.09 46.24 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 46.24 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 40.635 42.88 40.965 ;
      VIA 42.09 40.8 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 40.615 42.86 40.985 ;
      VIA 42.09 40.8 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 40.8 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 35.195 42.88 35.525 ;
      VIA 42.09 35.36 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 35.175 42.86 35.545 ;
      VIA 42.09 35.36 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 35.36 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 29.755 42.88 30.085 ;
      VIA 42.09 29.92 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 29.735 42.86 30.105 ;
      VIA 42.09 29.92 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 29.92 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 24.315 42.88 24.645 ;
      VIA 42.09 24.48 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 24.295 42.86 24.665 ;
      VIA 42.09 24.48 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 24.48 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 18.875 42.88 19.205 ;
      VIA 42.09 19.04 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 18.855 42.86 19.225 ;
      VIA 42.09 19.04 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 19.04 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 13.435 42.88 13.765 ;
      VIA 42.09 13.6 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 13.415 42.86 13.785 ;
      VIA 42.09 13.6 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 13.6 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 7.995 42.88 8.325 ;
      VIA 42.09 8.16 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 7.975 42.86 8.345 ;
      VIA 42.09 8.16 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 8.16 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 2.555 42.88 2.885 ;
      VIA 42.09 2.72 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 2.535 42.86 2.905 ;
      VIA 42.09 2.72 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 2.72 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 165.755 15.74 166.085 ;
      VIA 14.95 165.92 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 165.735 15.72 166.105 ;
      VIA 14.95 165.92 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 165.92 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 160.315 15.74 160.645 ;
      VIA 14.95 160.48 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 160.295 15.72 160.665 ;
      VIA 14.95 160.48 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 160.48 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 154.875 15.74 155.205 ;
      VIA 14.95 155.04 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 154.855 15.72 155.225 ;
      VIA 14.95 155.04 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 155.04 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 149.435 15.74 149.765 ;
      VIA 14.95 149.6 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 149.415 15.72 149.785 ;
      VIA 14.95 149.6 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 149.6 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 143.995 15.74 144.325 ;
      VIA 14.95 144.16 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 143.975 15.72 144.345 ;
      VIA 14.95 144.16 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 144.16 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 138.555 15.74 138.885 ;
      VIA 14.95 138.72 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 138.535 15.72 138.905 ;
      VIA 14.95 138.72 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 138.72 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 133.115 15.74 133.445 ;
      VIA 14.95 133.28 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 133.095 15.72 133.465 ;
      VIA 14.95 133.28 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 133.28 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 127.675 15.74 128.005 ;
      VIA 14.95 127.84 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 127.655 15.72 128.025 ;
      VIA 14.95 127.84 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 127.84 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 122.235 15.74 122.565 ;
      VIA 14.95 122.4 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 122.215 15.72 122.585 ;
      VIA 14.95 122.4 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 122.4 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 116.795 15.74 117.125 ;
      VIA 14.95 116.96 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 116.775 15.72 117.145 ;
      VIA 14.95 116.96 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 116.96 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 111.355 15.74 111.685 ;
      VIA 14.95 111.52 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 111.335 15.72 111.705 ;
      VIA 14.95 111.52 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 111.52 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 105.915 15.74 106.245 ;
      VIA 14.95 106.08 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 105.895 15.72 106.265 ;
      VIA 14.95 106.08 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 106.08 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 100.475 15.74 100.805 ;
      VIA 14.95 100.64 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 100.455 15.72 100.825 ;
      VIA 14.95 100.64 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 100.64 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 95.035 15.74 95.365 ;
      VIA 14.95 95.2 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 95.015 15.72 95.385 ;
      VIA 14.95 95.2 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 95.2 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 89.595 15.74 89.925 ;
      VIA 14.95 89.76 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 89.575 15.72 89.945 ;
      VIA 14.95 89.76 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 89.76 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 84.155 15.74 84.485 ;
      VIA 14.95 84.32 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 84.135 15.72 84.505 ;
      VIA 14.95 84.32 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 84.32 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 78.715 15.74 79.045 ;
      VIA 14.95 78.88 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 78.695 15.72 79.065 ;
      VIA 14.95 78.88 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 78.88 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 73.275 15.74 73.605 ;
      VIA 14.95 73.44 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 73.255 15.72 73.625 ;
      VIA 14.95 73.44 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 73.44 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 67.835 15.74 68.165 ;
      VIA 14.95 68 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 67.815 15.72 68.185 ;
      VIA 14.95 68 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 68 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 62.395 15.74 62.725 ;
      VIA 14.95 62.56 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 62.375 15.72 62.745 ;
      VIA 14.95 62.56 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 62.56 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 56.955 15.74 57.285 ;
      VIA 14.95 57.12 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 56.935 15.72 57.305 ;
      VIA 14.95 57.12 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 57.12 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 51.515 15.74 51.845 ;
      VIA 14.95 51.68 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 51.495 15.72 51.865 ;
      VIA 14.95 51.68 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 51.68 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 46.075 15.74 46.405 ;
      VIA 14.95 46.24 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 46.055 15.72 46.425 ;
      VIA 14.95 46.24 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 46.24 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 40.635 15.74 40.965 ;
      VIA 14.95 40.8 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 40.615 15.72 40.985 ;
      VIA 14.95 40.8 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 40.8 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 35.195 15.74 35.525 ;
      VIA 14.95 35.36 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 35.175 15.72 35.545 ;
      VIA 14.95 35.36 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 35.36 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 29.755 15.74 30.085 ;
      VIA 14.95 29.92 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 29.735 15.72 30.105 ;
      VIA 14.95 29.92 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 29.92 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 24.315 15.74 24.645 ;
      VIA 14.95 24.48 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 24.295 15.72 24.665 ;
      VIA 14.95 24.48 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 24.48 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 18.875 15.74 19.205 ;
      VIA 14.95 19.04 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 18.855 15.72 19.225 ;
      VIA 14.95 19.04 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 19.04 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 13.435 15.74 13.765 ;
      VIA 14.95 13.6 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 13.415 15.72 13.785 ;
      VIA 14.95 13.6 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 13.6 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 7.995 15.74 8.325 ;
      VIA 14.95 8.16 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 7.975 15.72 8.345 ;
      VIA 14.95 8.16 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 8.16 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 2.555 15.74 2.885 ;
      VIA 14.95 2.72 ibex_wb_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 2.535 15.72 2.905 ;
      VIA 14.95 2.72 ibex_wb_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 2.72 ibex_wb_stage_via2_3_1600_480_1_5_320_320 ;
    END
  END VSS
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  5.68 0 5.82 0.485 ;
    END
  END clk_i
  PIN en_wb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  49.84 0 49.98 0.485 ;
    END
  END en_wb_i
  PIN instr_done_wb_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  33.28 0 33.42 0.485 ;
    END
  END instr_done_wb_o
  PIN instr_is_compressed_id_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  48 0 48.14 0.485 ;
    END
  END instr_is_compressed_id_i
  PIN instr_perf_count_id_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  46.16 0 46.3 0.485 ;
    END
  END instr_perf_count_id_i
  PIN instr_type_wb_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  7.52 0 7.66 0.485 ;
    END
  END instr_type_wb_i[0]
  PIN instr_type_wb_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  9.36 0 9.5 0.485 ;
    END
  END instr_type_wb_i[1]
  PIN lsu_resp_err_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  44.32 0 44.46 0.485 ;
    END
  END lsu_resp_err_i
  PIN lsu_resp_valid_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  42.48 0 42.62 0.485 ;
    END
  END lsu_resp_valid_i
  PIN outstanding_load_wb_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 67.51 0.8 67.81 ;
    END
  END outstanding_load_wb_o
  PIN outstanding_store_wb_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 47.11 0.8 47.41 ;
    END
  END outstanding_store_wb_o
  PIN pc_id_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  11.2 0 11.34 0.485 ;
    END
  END pc_id_i[0]
  PIN pc_id_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  13.04 0 13.18 0.485 ;
    END
  END pc_id_i[10]
  PIN pc_id_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  14.88 0 15.02 0.485 ;
    END
  END pc_id_i[11]
  PIN pc_id_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  16.72 0 16.86 0.485 ;
    END
  END pc_id_i[12]
  PIN pc_id_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  18.56 0 18.7 0.485 ;
    END
  END pc_id_i[13]
  PIN pc_id_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  20.4 0 20.54 0.485 ;
    END
  END pc_id_i[14]
  PIN pc_id_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  22.24 0 22.38 0.485 ;
    END
  END pc_id_i[15]
  PIN pc_id_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  24.08 0 24.22 0.485 ;
    END
  END pc_id_i[16]
  PIN pc_id_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  25.92 0 26.06 0.485 ;
    END
  END pc_id_i[17]
  PIN pc_id_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  27.76 0 27.9 0.485 ;
    END
  END pc_id_i[18]
  PIN pc_id_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  29.6 0 29.74 0.485 ;
    END
  END pc_id_i[19]
  PIN pc_id_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  31.44 0 31.58 0.485 ;
    END
  END pc_id_i[1]
  PIN pc_id_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  2 0 2.14 0.485 ;
    END
  END pc_id_i[20]
  PIN pc_id_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  35.12 0 35.26 0.485 ;
    END
  END pc_id_i[21]
  PIN pc_id_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  36.96 0 37.1 0.485 ;
    END
  END pc_id_i[22]
  PIN pc_id_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  38.8 0 38.94 0.485 ;
    END
  END pc_id_i[23]
  PIN pc_id_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  40.64 0 40.78 0.485 ;
    END
  END pc_id_i[24]
  PIN pc_id_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  53.52 0 53.66 0.485 ;
    END
  END pc_id_i[25]
  PIN pc_id_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  51.68 0 51.82 0.485 ;
    END
  END pc_id_i[26]
  PIN pc_id_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  55.36 0 55.5 0.485 ;
    END
  END pc_id_i[27]
  PIN pc_id_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  3.84 0 3.98 0.485 ;
    END
  END pc_id_i[28]
  PIN pc_id_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 155.23 58.02 155.53 ;
    END
  END pc_id_i[29]
  PIN pc_id_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 161.35 58.02 161.65 ;
    END
  END pc_id_i[2]
  PIN pc_id_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 4.27 58.02 4.57 ;
    END
  END pc_id_i[30]
  PIN pc_id_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 167.47 58.02 167.77 ;
    END
  END pc_id_i[31]
  PIN pc_id_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 20.59 58.02 20.89 ;
    END
  END pc_id_i[3]
  PIN pc_id_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 163.39 58.02 163.69 ;
    END
  END pc_id_i[4]
  PIN pc_id_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 18.55 58.02 18.85 ;
    END
  END pc_id_i[5]
  PIN pc_id_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 157.27 58.02 157.57 ;
    END
  END pc_id_i[6]
  PIN pc_id_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 2.23 58.02 2.53 ;
    END
  END pc_id_i[7]
  PIN pc_id_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 165.43 58.02 165.73 ;
    END
  END pc_id_i[8]
  PIN pc_id_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 159.31 58.02 159.61 ;
    END
  END pc_id_i[9]
  PIN pc_wb_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 34.87 0.8 35.17 ;
    END
  END pc_wb_o[0]
  PIN pc_wb_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 32.83 0.8 33.13 ;
    END
  END pc_wb_o[10]
  PIN pc_wb_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 18.55 0.8 18.85 ;
    END
  END pc_wb_o[11]
  PIN pc_wb_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 40.99 58.02 41.29 ;
    END
  END pc_wb_o[12]
  PIN pc_wb_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 22.63 58.02 22.93 ;
    END
  END pc_wb_o[13]
  PIN pc_wb_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 91.99 58.02 92.29 ;
    END
  END pc_wb_o[14]
  PIN pc_wb_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 20.59 0.8 20.89 ;
    END
  END pc_wb_o[15]
  PIN pc_wb_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 47.11 58.02 47.41 ;
    END
  END pc_wb_o[16]
  PIN pc_wb_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 36.91 0.8 37.21 ;
    END
  END pc_wb_o[17]
  PIN pc_wb_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 51.19 58.02 51.49 ;
    END
  END pc_wb_o[18]
  PIN pc_wb_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 73.63 0.8 73.93 ;
    END
  END pc_wb_o[19]
  PIN pc_wb_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 71.59 58.02 71.89 ;
    END
  END pc_wb_o[1]
  PIN pc_wb_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 30.79 58.02 31.09 ;
    END
  END pc_wb_o[20]
  PIN pc_wb_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 30.79 0.8 31.09 ;
    END
  END pc_wb_o[21]
  PIN pc_wb_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 55.27 58.02 55.57 ;
    END
  END pc_wb_o[22]
  PIN pc_wb_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 77.71 0.8 78.01 ;
    END
  END pc_wb_o[23]
  PIN pc_wb_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 24.67 0.8 24.97 ;
    END
  END pc_wb_o[24]
  PIN pc_wb_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 87.91 58.02 88.21 ;
    END
  END pc_wb_o[25]
  PIN pc_wb_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 65.47 58.02 65.77 ;
    END
  END pc_wb_o[26]
  PIN pc_wb_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 79.75 58.02 80.05 ;
    END
  END pc_wb_o[27]
  PIN pc_wb_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 57.31 58.02 57.61 ;
    END
  END pc_wb_o[28]
  PIN pc_wb_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 45.07 0.8 45.37 ;
    END
  END pc_wb_o[29]
  PIN pc_wb_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 59.35 58.02 59.65 ;
    END
  END pc_wb_o[2]
  PIN pc_wb_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 26.71 0.8 27.01 ;
    END
  END pc_wb_o[30]
  PIN pc_wb_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 71.59 0.8 71.89 ;
    END
  END pc_wb_o[31]
  PIN pc_wb_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 65.47 0.8 65.77 ;
    END
  END pc_wb_o[3]
  PIN pc_wb_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 79.75 0.8 80.05 ;
    END
  END pc_wb_o[4]
  PIN pc_wb_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 75.67 58.02 75.97 ;
    END
  END pc_wb_o[5]
  PIN pc_wb_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 40.99 0.8 41.29 ;
    END
  END pc_wb_o[6]
  PIN pc_wb_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 67.51 58.02 67.81 ;
    END
  END pc_wb_o[7]
  PIN pc_wb_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 61.39 58.02 61.69 ;
    END
  END pc_wb_o[8]
  PIN pc_wb_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 49.15 58.02 49.45 ;
    END
  END pc_wb_o[9]
  PIN perf_instr_ret_compressed_wb_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 16.51 58.02 16.81 ;
    END
  END perf_instr_ret_compressed_wb_o
  PIN perf_instr_ret_wb_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 14.47 58.02 14.77 ;
    END
  END perf_instr_ret_wb_o
  PIN ready_wb_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  2 169.58 2.14 170.065 ;
    END
  END ready_wb_o
  PIN rf_waddr_id_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  3.84 169.58 3.98 170.065 ;
    END
  END rf_waddr_id_i[0]
  PIN rf_waddr_id_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 8.35 0.8 8.65 ;
    END
  END rf_waddr_id_i[1]
  PIN rf_waddr_id_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 10.39 58.02 10.69 ;
    END
  END rf_waddr_id_i[2]
  PIN rf_waddr_id_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 10.39 0.8 10.69 ;
    END
  END rf_waddr_id_i[3]
  PIN rf_waddr_id_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 6.31 58.02 6.61 ;
    END
  END rf_waddr_id_i[4]
  PIN rf_waddr_wb_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  7.52 169.58 7.66 170.065 ;
    END
  END rf_waddr_wb_o[0]
  PIN rf_waddr_wb_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 14.47 0.8 14.77 ;
    END
  END rf_waddr_wb_o[1]
  PIN rf_waddr_wb_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 12.43 58.02 12.73 ;
    END
  END rf_waddr_wb_o[2]
  PIN rf_waddr_wb_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 12.43 0.8 12.73 ;
    END
  END rf_waddr_wb_o[3]
  PIN rf_waddr_wb_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 8.35 58.02 8.65 ;
    END
  END rf_waddr_wb_o[4]
  PIN rf_wdata_fwd_wb_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 53.23 58.02 53.53 ;
    END
  END rf_wdata_fwd_wb_o[0]
  PIN rf_wdata_fwd_wb_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 81.79 58.02 82.09 ;
    END
  END rf_wdata_fwd_wb_o[10]
  PIN rf_wdata_fwd_wb_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 55.27 0.8 55.57 ;
    END
  END rf_wdata_fwd_wb_o[11]
  PIN rf_wdata_fwd_wb_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 63.43 0.8 63.73 ;
    END
  END rf_wdata_fwd_wb_o[12]
  PIN rf_wdata_fwd_wb_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 77.71 58.02 78.01 ;
    END
  END rf_wdata_fwd_wb_o[13]
  PIN rf_wdata_fwd_wb_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 75.67 0.8 75.97 ;
    END
  END rf_wdata_fwd_wb_o[14]
  PIN rf_wdata_fwd_wb_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 26.71 58.02 27.01 ;
    END
  END rf_wdata_fwd_wb_o[15]
  PIN rf_wdata_fwd_wb_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 38.95 58.02 39.25 ;
    END
  END rf_wdata_fwd_wb_o[16]
  PIN rf_wdata_fwd_wb_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 85.87 58.02 86.17 ;
    END
  END rf_wdata_fwd_wb_o[17]
  PIN rf_wdata_fwd_wb_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 43.03 58.02 43.33 ;
    END
  END rf_wdata_fwd_wb_o[18]
  PIN rf_wdata_fwd_wb_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 22.63 0.8 22.93 ;
    END
  END rf_wdata_fwd_wb_o[19]
  PIN rf_wdata_fwd_wb_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 34.87 58.02 35.17 ;
    END
  END rf_wdata_fwd_wb_o[1]
  PIN rf_wdata_fwd_wb_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 51.19 0.8 51.49 ;
    END
  END rf_wdata_fwd_wb_o[20]
  PIN rf_wdata_fwd_wb_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 32.83 58.02 33.13 ;
    END
  END rf_wdata_fwd_wb_o[21]
  PIN rf_wdata_fwd_wb_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 59.35 0.8 59.65 ;
    END
  END rf_wdata_fwd_wb_o[22]
  PIN rf_wdata_fwd_wb_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 61.39 0.8 61.69 ;
    END
  END rf_wdata_fwd_wb_o[23]
  PIN rf_wdata_fwd_wb_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 69.55 0.8 69.85 ;
    END
  END rf_wdata_fwd_wb_o[24]
  PIN rf_wdata_fwd_wb_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 89.95 58.02 90.25 ;
    END
  END rf_wdata_fwd_wb_o[25]
  PIN rf_wdata_fwd_wb_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 36.91 58.02 37.21 ;
    END
  END rf_wdata_fwd_wb_o[26]
  PIN rf_wdata_fwd_wb_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 43.03 0.8 43.33 ;
    END
  END rf_wdata_fwd_wb_o[27]
  PIN rf_wdata_fwd_wb_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 28.75 0.8 29.05 ;
    END
  END rf_wdata_fwd_wb_o[28]
  PIN rf_wdata_fwd_wb_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 45.07 58.02 45.37 ;
    END
  END rf_wdata_fwd_wb_o[29]
  PIN rf_wdata_fwd_wb_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 69.55 58.02 69.85 ;
    END
  END rf_wdata_fwd_wb_o[2]
  PIN rf_wdata_fwd_wb_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 83.83 58.02 84.13 ;
    END
  END rf_wdata_fwd_wb_o[30]
  PIN rf_wdata_fwd_wb_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 63.43 58.02 63.73 ;
    END
  END rf_wdata_fwd_wb_o[31]
  PIN rf_wdata_fwd_wb_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 53.23 0.8 53.53 ;
    END
  END rf_wdata_fwd_wb_o[3]
  PIN rf_wdata_fwd_wb_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 81.79 0.8 82.09 ;
    END
  END rf_wdata_fwd_wb_o[4]
  PIN rf_wdata_fwd_wb_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 57.31 0.8 57.61 ;
    END
  END rf_wdata_fwd_wb_o[5]
  PIN rf_wdata_fwd_wb_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 73.63 58.02 73.93 ;
    END
  END rf_wdata_fwd_wb_o[6]
  PIN rf_wdata_fwd_wb_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 24.67 58.02 24.97 ;
    END
  END rf_wdata_fwd_wb_o[7]
  PIN rf_wdata_fwd_wb_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 28.75 58.02 29.05 ;
    END
  END rf_wdata_fwd_wb_o[8]
  PIN rf_wdata_fwd_wb_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 38.95 0.8 39.25 ;
    END
  END rf_wdata_fwd_wb_o[9]
  PIN rf_wdata_id_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 157.27 0.8 157.57 ;
    END
  END rf_wdata_id_i[0]
  PIN rf_wdata_id_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 120.55 0.8 120.85 ;
    END
  END rf_wdata_id_i[10]
  PIN rf_wdata_id_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 85.87 0.8 86.17 ;
    END
  END rf_wdata_id_i[11]
  PIN rf_wdata_id_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 91.99 0.8 92.29 ;
    END
  END rf_wdata_id_i[12]
  PIN rf_wdata_id_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 100.15 0.8 100.45 ;
    END
  END rf_wdata_id_i[13]
  PIN rf_wdata_id_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 134.83 0.8 135.13 ;
    END
  END rf_wdata_id_i[14]
  PIN rf_wdata_id_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 96.07 0.8 96.37 ;
    END
  END rf_wdata_id_i[15]
  PIN rf_wdata_id_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 124.63 0.8 124.93 ;
    END
  END rf_wdata_id_i[16]
  PIN rf_wdata_id_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 110.35 0.8 110.65 ;
    END
  END rf_wdata_id_i[17]
  PIN rf_wdata_id_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 153.19 58.02 153.49 ;
    END
  END rf_wdata_id_i[18]
  PIN rf_wdata_id_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 147.07 58.02 147.37 ;
    END
  END rf_wdata_id_i[19]
  PIN rf_wdata_id_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 110.35 58.02 110.65 ;
    END
  END rf_wdata_id_i[1]
  PIN rf_wdata_id_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 149.11 58.02 149.41 ;
    END
  END rf_wdata_id_i[20]
  PIN rf_wdata_id_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 145.03 58.02 145.33 ;
    END
  END rf_wdata_id_i[21]
  PIN rf_wdata_id_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 98.11 58.02 98.41 ;
    END
  END rf_wdata_id_i[22]
  PIN rf_wdata_id_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 112.39 58.02 112.69 ;
    END
  END rf_wdata_id_i[23]
  PIN rf_wdata_id_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 106.27 58.02 106.57 ;
    END
  END rf_wdata_id_i[24]
  PIN rf_wdata_id_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 138.91 58.02 139.21 ;
    END
  END rf_wdata_id_i[25]
  PIN rf_wdata_id_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 116.47 58.02 116.77 ;
    END
  END rf_wdata_id_i[26]
  PIN rf_wdata_id_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  40.64 169.58 40.78 170.065 ;
    END
  END rf_wdata_id_i[27]
  PIN rf_wdata_id_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  9.36 169.58 9.5 170.065 ;
    END
  END rf_wdata_id_i[28]
  PIN rf_wdata_id_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  48 169.58 48.14 170.065 ;
    END
  END rf_wdata_id_i[29]
  PIN rf_wdata_id_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  51.68 169.58 51.82 170.065 ;
    END
  END rf_wdata_id_i[2]
  PIN rf_wdata_id_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  55.36 169.58 55.5 170.065 ;
    END
  END rf_wdata_id_i[30]
  PIN rf_wdata_id_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  53.52 169.58 53.66 170.065 ;
    END
  END rf_wdata_id_i[31]
  PIN rf_wdata_id_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  35.12 169.58 35.26 170.065 ;
    END
  END rf_wdata_id_i[3]
  PIN rf_wdata_id_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  31.44 169.58 31.58 170.065 ;
    END
  END rf_wdata_id_i[4]
  PIN rf_wdata_id_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  16.72 169.58 16.86 170.065 ;
    END
  END rf_wdata_id_i[5]
  PIN rf_wdata_id_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  29.6 169.58 29.74 170.065 ;
    END
  END rf_wdata_id_i[6]
  PIN rf_wdata_id_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  14.88 169.58 15.02 170.065 ;
    END
  END rf_wdata_id_i[7]
  PIN rf_wdata_id_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  11.2 169.58 11.34 170.065 ;
    END
  END rf_wdata_id_i[8]
  PIN rf_wdata_id_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  24.08 169.58 24.22 170.065 ;
    END
  END rf_wdata_id_i[9]
  PIN rf_wdata_lsu_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 116.47 0.8 116.77 ;
    END
  END rf_wdata_lsu_i[0]
  PIN rf_wdata_lsu_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 112.39 0.8 112.69 ;
    END
  END rf_wdata_lsu_i[10]
  PIN rf_wdata_lsu_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 106.27 0.8 106.57 ;
    END
  END rf_wdata_lsu_i[11]
  PIN rf_wdata_lsu_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 94.03 0.8 94.33 ;
    END
  END rf_wdata_lsu_i[12]
  PIN rf_wdata_lsu_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 89.95 0.8 90.25 ;
    END
  END rf_wdata_lsu_i[13]
  PIN rf_wdata_lsu_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 126.67 0.8 126.97 ;
    END
  END rf_wdata_lsu_i[14]
  PIN rf_wdata_lsu_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 104.23 0.8 104.53 ;
    END
  END rf_wdata_lsu_i[15]
  PIN rf_wdata_lsu_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 128.71 0.8 129.01 ;
    END
  END rf_wdata_lsu_i[16]
  PIN rf_wdata_lsu_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 118.51 0.8 118.81 ;
    END
  END rf_wdata_lsu_i[17]
  PIN rf_wdata_lsu_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 122.59 58.02 122.89 ;
    END
  END rf_wdata_lsu_i[18]
  PIN rf_wdata_lsu_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 124.63 58.02 124.93 ;
    END
  END rf_wdata_lsu_i[19]
  PIN rf_wdata_lsu_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 102.19 58.02 102.49 ;
    END
  END rf_wdata_lsu_i[1]
  PIN rf_wdata_lsu_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 134.83 58.02 135.13 ;
    END
  END rf_wdata_lsu_i[20]
  PIN rf_wdata_lsu_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 142.99 58.02 143.29 ;
    END
  END rf_wdata_lsu_i[21]
  PIN rf_wdata_lsu_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 94.03 58.02 94.33 ;
    END
  END rf_wdata_lsu_i[22]
  PIN rf_wdata_lsu_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 114.43 58.02 114.73 ;
    END
  END rf_wdata_lsu_i[23]
  PIN rf_wdata_lsu_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 96.07 58.02 96.37 ;
    END
  END rf_wdata_lsu_i[24]
  PIN rf_wdata_lsu_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 136.87 58.02 137.17 ;
    END
  END rf_wdata_lsu_i[25]
  PIN rf_wdata_lsu_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 126.67 58.02 126.97 ;
    END
  END rf_wdata_lsu_i[26]
  PIN rf_wdata_lsu_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  38.8 169.58 38.94 170.065 ;
    END
  END rf_wdata_lsu_i[27]
  PIN rf_wdata_lsu_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  20.4 169.58 20.54 170.065 ;
    END
  END rf_wdata_lsu_i[28]
  PIN rf_wdata_lsu_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  44.32 169.58 44.46 170.065 ;
    END
  END rf_wdata_lsu_i[29]
  PIN rf_wdata_lsu_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  49.84 169.58 49.98 170.065 ;
    END
  END rf_wdata_lsu_i[2]
  PIN rf_wdata_lsu_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  42.48 169.58 42.62 170.065 ;
    END
  END rf_wdata_lsu_i[30]
  PIN rf_wdata_lsu_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  46.16 169.58 46.3 170.065 ;
    END
  END rf_wdata_lsu_i[31]
  PIN rf_wdata_lsu_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  36.96 169.58 37.1 170.065 ;
    END
  END rf_wdata_lsu_i[3]
  PIN rf_wdata_lsu_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  33.28 169.58 33.42 170.065 ;
    END
  END rf_wdata_lsu_i[4]
  PIN rf_wdata_lsu_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  25.92 169.58 26.06 170.065 ;
    END
  END rf_wdata_lsu_i[5]
  PIN rf_wdata_lsu_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  27.76 169.58 27.9 170.065 ;
    END
  END rf_wdata_lsu_i[6]
  PIN rf_wdata_lsu_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  18.56 169.58 18.7 170.065 ;
    END
  END rf_wdata_lsu_i[7]
  PIN rf_wdata_lsu_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  13.04 169.58 13.18 170.065 ;
    END
  END rf_wdata_lsu_i[8]
  PIN rf_wdata_lsu_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  5.68 169.58 5.82 170.065 ;
    END
  END rf_wdata_lsu_i[9]
  PIN rf_wdata_wb_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  22.24 169.58 22.38 170.065 ;
    END
  END rf_wdata_wb_o[0]
  PIN rf_wdata_wb_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 114.43 0.8 114.73 ;
    END
  END rf_wdata_wb_o[10]
  PIN rf_wdata_wb_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 83.83 0.8 84.13 ;
    END
  END rf_wdata_wb_o[11]
  PIN rf_wdata_wb_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 98.11 0.8 98.41 ;
    END
  END rf_wdata_wb_o[12]
  PIN rf_wdata_wb_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 87.91 0.8 88.21 ;
    END
  END rf_wdata_wb_o[13]
  PIN rf_wdata_wb_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 130.75 0.8 131.05 ;
    END
  END rf_wdata_wb_o[14]
  PIN rf_wdata_wb_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 102.19 0.8 102.49 ;
    END
  END rf_wdata_wb_o[15]
  PIN rf_wdata_wb_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 122.59 0.8 122.89 ;
    END
  END rf_wdata_wb_o[16]
  PIN rf_wdata_wb_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 108.31 0.8 108.61 ;
    END
  END rf_wdata_wb_o[17]
  PIN rf_wdata_wb_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 120.55 58.02 120.85 ;
    END
  END rf_wdata_wb_o[18]
  PIN rf_wdata_wb_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 151.15 58.02 151.45 ;
    END
  END rf_wdata_wb_o[19]
  PIN rf_wdata_wb_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 104.23 58.02 104.53 ;
    END
  END rf_wdata_wb_o[1]
  PIN rf_wdata_wb_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 130.75 58.02 131.05 ;
    END
  END rf_wdata_wb_o[20]
  PIN rf_wdata_wb_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 132.79 58.02 133.09 ;
    END
  END rf_wdata_wb_o[21]
  PIN rf_wdata_wb_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 108.31 58.02 108.61 ;
    END
  END rf_wdata_wb_o[22]
  PIN rf_wdata_wb_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 118.51 58.02 118.81 ;
    END
  END rf_wdata_wb_o[23]
  PIN rf_wdata_wb_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 100.15 58.02 100.45 ;
    END
  END rf_wdata_wb_o[24]
  PIN rf_wdata_wb_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 140.95 58.02 141.25 ;
    END
  END rf_wdata_wb_o[25]
  PIN rf_wdata_wb_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  57.22 128.71 58.02 129.01 ;
    END
  END rf_wdata_wb_o[26]
  PIN rf_wdata_wb_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 149.11 0.8 149.41 ;
    END
  END rf_wdata_wb_o[27]
  PIN rf_wdata_wb_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 155.23 0.8 155.53 ;
    END
  END rf_wdata_wb_o[28]
  PIN rf_wdata_wb_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 167.47 0.8 167.77 ;
    END
  END rf_wdata_wb_o[29]
  PIN rf_wdata_wb_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 153.19 0.8 153.49 ;
    END
  END rf_wdata_wb_o[2]
  PIN rf_wdata_wb_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 142.99 0.8 143.29 ;
    END
  END rf_wdata_wb_o[30]
  PIN rf_wdata_wb_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 161.35 0.8 161.65 ;
    END
  END rf_wdata_wb_o[31]
  PIN rf_wdata_wb_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 140.95 0.8 141.25 ;
    END
  END rf_wdata_wb_o[3]
  PIN rf_wdata_wb_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 163.39 0.8 163.69 ;
    END
  END rf_wdata_wb_o[4]
  PIN rf_wdata_wb_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 165.43 0.8 165.73 ;
    END
  END rf_wdata_wb_o[5]
  PIN rf_wdata_wb_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 159.31 0.8 159.61 ;
    END
  END rf_wdata_wb_o[6]
  PIN rf_wdata_wb_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 138.91 0.8 139.21 ;
    END
  END rf_wdata_wb_o[7]
  PIN rf_wdata_wb_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 145.03 0.8 145.33 ;
    END
  END rf_wdata_wb_o[8]
  PIN rf_wdata_wb_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 147.07 0.8 147.37 ;
    END
  END rf_wdata_wb_o[9]
  PIN rf_we_id_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 151.15 0.8 151.45 ;
    END
  END rf_we_id_i
  PIN rf_we_lsu_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 136.87 0.8 137.17 ;
    END
  END rf_we_lsu_i
  PIN rf_we_wb_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 132.79 0.8 133.09 ;
    END
  END rf_we_wb_o
  PIN rf_write_wb_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 49.15 0.8 49.45 ;
    END
  END rf_write_wb_o
  PIN rst_ni
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 16.51 0.8 16.81 ;
    END
  END rst_ni
  OBS
    LAYER nwell ;
     RECT  0 0 58.02 170.065 ;
    LAYER pwell ;
     RECT  0 0 58.02 170.065 ;
    LAYER li1 ;
     RECT  0 0 58.02 170.065 ;
    LAYER met1 ;
     RECT  0 0 58.02 170.065 ;
    LAYER met2 ;
     RECT  0 0 58.02 170.065 ;
    LAYER met3 ;
     RECT  0 0 58.02 170.065 ;
    LAYER met4 ;
     RECT  0 0 58.02 170.065 ;
    LAYER met5 ;
     RECT  0 0 58.02 170.065 ;
  END
END ibex_wb_stage
END LIBRARY
