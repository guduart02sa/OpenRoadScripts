module ibex_if_stage (clk_i,
    csr_mtvec_init_o,
    dummy_instr_en_i,
    dummy_instr_id_o,
    dummy_instr_seed_en_i,
    icache_enable_i,
    icache_inval_i,
    id_in_ready_i,
    if_busy_o,
    illegal_c_insn_id_o,
    instr_bp_taken_o,
    instr_err_i,
    instr_fetch_err_o,
    instr_fetch_err_plus2_o,
    instr_gnt_i,
    instr_is_compressed_id_o,
    instr_new_id_o,
    instr_pmp_err_i,
    instr_req_o,
    instr_rvalid_i,
    instr_valid_clear_i,
    instr_valid_id_o,
    nt_branch_mispredict_i,
    pc_mismatch_alert_o,
    pc_set_i,
    pc_set_spec_i,
    req_i,
    rst_ni,
    boot_addr_i,
    branch_target_ex_i,
    csr_depc_i,
    csr_mepc_i,
    csr_mtvec_i,
    dummy_instr_mask_i,
    dummy_instr_seed_i,
    exc_cause,
    exc_pc_mux_i,
    instr_addr_o,
    instr_rdata_alu_id_o,
    instr_rdata_c_id_o,
    instr_rdata_i,
    instr_rdata_id_o,
    pc_id_o,
    pc_if_o,
    pc_mux_i);
 input clk_i;
 output csr_mtvec_init_o;
 input dummy_instr_en_i;
 output dummy_instr_id_o;
 input dummy_instr_seed_en_i;
 input icache_enable_i;
 input icache_inval_i;
 input id_in_ready_i;
 output if_busy_o;
 output illegal_c_insn_id_o;
 output instr_bp_taken_o;
 input instr_err_i;
 output instr_fetch_err_o;
 output instr_fetch_err_plus2_o;
 input instr_gnt_i;
 output instr_is_compressed_id_o;
 output instr_new_id_o;
 input instr_pmp_err_i;
 output instr_req_o;
 input instr_rvalid_i;
 input instr_valid_clear_i;
 output instr_valid_id_o;
 input nt_branch_mispredict_i;
 output pc_mismatch_alert_o;
 input pc_set_i;
 input pc_set_spec_i;
 input req_i;
 input rst_ni;
 input [31:0] boot_addr_i;
 input [31:0] branch_target_ex_i;
 input [31:0] csr_depc_i;
 input [31:0] csr_mepc_i;
 input [31:0] csr_mtvec_i;
 input [2:0] dummy_instr_mask_i;
 input [31:0] dummy_instr_seed_i;
 input [5:0] exc_cause;
 input [1:0] exc_pc_mux_i;
 output [31:0] instr_addr_o;
 output [31:0] instr_rdata_alu_id_o;
 output [15:0] instr_rdata_c_id_o;
 input [31:0] instr_rdata_i;
 output [31:0] instr_rdata_id_o;
 output [31:0] pc_id_o;
 output [31:0] pc_if_o;
 input [2:0] pc_mux_i;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire clknet_leaf_0_clk_i;
 wire \compressed_decoder_i.illegal_instr_o ;
 wire \compressed_decoder_i.instr_i[0] ;
 wire \compressed_decoder_i.instr_i[10] ;
 wire \compressed_decoder_i.instr_i[11] ;
 wire \compressed_decoder_i.instr_i[12] ;
 wire \compressed_decoder_i.instr_i[13] ;
 wire \compressed_decoder_i.instr_i[14] ;
 wire \compressed_decoder_i.instr_i[15] ;
 wire \compressed_decoder_i.instr_i[1] ;
 wire \compressed_decoder_i.instr_i[2] ;
 wire \compressed_decoder_i.instr_i[3] ;
 wire \compressed_decoder_i.instr_i[4] ;
 wire \compressed_decoder_i.instr_i[5] ;
 wire \compressed_decoder_i.instr_i[6] ;
 wire \compressed_decoder_i.instr_i[7] ;
 wire \compressed_decoder_i.instr_i[8] ;
 wire \compressed_decoder_i.instr_i[9] ;
 wire \compressed_decoder_i.instr_o[0] ;
 wire \compressed_decoder_i.instr_o[10] ;
 wire \compressed_decoder_i.instr_o[11] ;
 wire \compressed_decoder_i.instr_o[12] ;
 wire \compressed_decoder_i.instr_o[13] ;
 wire \compressed_decoder_i.instr_o[14] ;
 wire \compressed_decoder_i.instr_o[15] ;
 wire \compressed_decoder_i.instr_o[16] ;
 wire \compressed_decoder_i.instr_o[17] ;
 wire \compressed_decoder_i.instr_o[18] ;
 wire \compressed_decoder_i.instr_o[19] ;
 wire \compressed_decoder_i.instr_o[1] ;
 wire \compressed_decoder_i.instr_o[20] ;
 wire \compressed_decoder_i.instr_o[21] ;
 wire \compressed_decoder_i.instr_o[22] ;
 wire \compressed_decoder_i.instr_o[23] ;
 wire \compressed_decoder_i.instr_o[24] ;
 wire \compressed_decoder_i.instr_o[25] ;
 wire \compressed_decoder_i.instr_o[26] ;
 wire \compressed_decoder_i.instr_o[27] ;
 wire \compressed_decoder_i.instr_o[28] ;
 wire \compressed_decoder_i.instr_o[29] ;
 wire \compressed_decoder_i.instr_o[2] ;
 wire \compressed_decoder_i.instr_o[30] ;
 wire \compressed_decoder_i.instr_o[31] ;
 wire \compressed_decoder_i.instr_o[3] ;
 wire \compressed_decoder_i.instr_o[4] ;
 wire \compressed_decoder_i.instr_o[5] ;
 wire \compressed_decoder_i.instr_o[6] ;
 wire \compressed_decoder_i.instr_o[7] ;
 wire \compressed_decoder_i.instr_o[8] ;
 wire \compressed_decoder_i.instr_o[9] ;
 wire \compressed_decoder_i.is_compressed_o ;
 wire net198;
 wire fetch_err;
 wire \gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[1] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[0] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[1] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.discard_req_d ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.discard_req_q ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[10] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[11] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[12] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[13] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[14] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[15] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[16] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[17] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[18] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[19] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[20] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[21] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[22] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[23] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[24] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[25] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[26] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[27] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[28] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[29] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[2] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[30] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[31] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[3] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[4] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[5] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[6] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[7] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[8] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[9] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[10] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[11] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[12] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[13] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[14] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[15] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[16] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[17] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[18] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[19] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[20] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[21] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[22] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[23] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[24] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[25] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[26] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[27] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[28] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[29] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[2] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[30] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[31] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[3] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[4] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[5] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[6] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[7] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[8] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[9] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[1] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[2] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_d[0] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_d[1] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_d[2] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[0] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[2] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[10] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[11] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[12] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[13] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[14] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[15] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[16] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[17] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[18] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[19] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[1] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[20] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[21] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[22] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[23] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[24] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[25] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[26] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[27] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[28] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[29] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[2] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[30] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[31] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[3] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[4] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[5] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[6] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[7] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[8] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[9] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_en ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[0] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[10] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[11] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[12] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[13] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[14] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[15] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[16] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[17] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[18] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[19] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[1] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[20] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[21] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[22] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[23] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[24] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[25] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[26] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[27] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[28] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[29] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[2] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[30] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[31] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[32] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[33] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[34] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[35] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[36] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[37] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[38] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[39] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[3] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[40] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[41] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[42] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[43] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[44] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[45] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[46] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[47] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[48] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[49] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[4] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[50] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[51] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[52] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[53] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[54] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[55] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[56] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[57] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[58] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[59] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[5] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[60] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[61] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[62] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[63] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[6] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[7] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[8] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[9] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[0] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[10] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[11] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[12] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[13] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[14] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[15] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[16] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[17] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[18] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[19] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[1] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[20] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[21] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[22] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[23] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[24] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[25] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[26] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[27] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[28] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[29] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[2] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[30] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[31] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[32] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[33] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[34] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[35] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[36] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[37] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[38] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[39] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[3] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[40] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[41] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[42] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[43] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[44] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[45] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[46] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[47] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[48] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[49] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[4] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[50] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[51] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[52] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[53] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[54] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[55] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[56] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[57] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[58] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[59] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[5] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[60] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[61] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[62] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[63] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[64] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[65] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[66] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[67] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[68] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[69] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[6] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[70] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[71] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[72] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[73] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[74] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[75] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[76] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[77] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[78] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[79] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[7] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[80] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[81] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[82] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[83] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[84] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[85] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[86] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[87] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[88] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[89] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[8] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[90] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[91] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[92] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[93] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[94] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[95] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[9] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[0] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[1] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[2] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[0] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[1] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.rdata_pmp_err_q[0] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.rdata_pmp_err_q[1] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.rdata_pmp_err_s[0] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.rdata_pmp_err_s[1] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[10] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[11] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[12] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[13] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[14] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[15] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[16] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[17] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[18] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[19] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[20] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[21] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[22] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[23] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[24] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[25] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[26] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[27] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[28] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[29] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[2] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[30] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[31] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[3] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[4] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[5] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[6] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[7] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[8] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[9] ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.valid_req_d ;
 wire \gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ;
 wire net199;
 wire if_id_pipe_reg_we;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire instr_valid_id_d;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire clknet_leaf_1_clk_i;
 wire clknet_leaf_2_clk_i;
 wire clknet_leaf_3_clk_i;
 wire clknet_leaf_4_clk_i;
 wire clknet_leaf_5_clk_i;
 wire clknet_leaf_6_clk_i;
 wire clknet_leaf_7_clk_i;
 wire clknet_leaf_8_clk_i;
 wire clknet_leaf_9_clk_i;
 wire clknet_leaf_10_clk_i;
 wire clknet_leaf_11_clk_i;
 wire clknet_leaf_12_clk_i;
 wire clknet_leaf_13_clk_i;
 wire clknet_leaf_14_clk_i;
 wire clknet_leaf_15_clk_i;
 wire clknet_leaf_16_clk_i;
 wire clknet_leaf_17_clk_i;
 wire clknet_leaf_18_clk_i;
 wire clknet_leaf_19_clk_i;
 wire clknet_leaf_20_clk_i;
 wire clknet_leaf_21_clk_i;
 wire clknet_leaf_22_clk_i;
 wire clknet_leaf_23_clk_i;
 wire clknet_leaf_24_clk_i;
 wire clknet_leaf_25_clk_i;
 wire clknet_leaf_26_clk_i;
 wire clknet_leaf_27_clk_i;
 wire clknet_leaf_28_clk_i;
 wire clknet_leaf_29_clk_i;
 wire clknet_leaf_30_clk_i;
 wire clknet_leaf_31_clk_i;
 wire clknet_leaf_32_clk_i;
 wire clknet_leaf_33_clk_i;
 wire clknet_leaf_34_clk_i;
 wire clknet_0_clk_i;
 wire clknet_2_0__leaf_clk_i;
 wire clknet_2_1__leaf_clk_i;
 wire clknet_2_2__leaf_clk_i;
 wire clknet_2_3__leaf_clk_i;

 sky130_fd_sc_hd__buf_4 _1070_ (.A(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .X(_0745_));
 sky130_fd_sc_hd__clkbuf_8 _1071_ (.A(_0745_),
    .X(_0746_));
 sky130_fd_sc_hd__buf_6 _1072_ (.A(_0746_),
    .X(_0747_));
 sky130_fd_sc_hd__mux2_2 _1073_ (.A0(net166),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[17] ),
    .S(_0747_),
    .X(_0748_));
 sky130_fd_sc_hd__mux2_1 _1074_ (.A0(net169),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[1] ),
    .S(_0747_),
    .X(_0749_));
 sky130_fd_sc_hd__inv_6 _1075_ (.A(net358),
    .Y(_0750_));
 sky130_fd_sc_hd__buf_8 _1076_ (.A(_0750_),
    .X(_0751_));
 sky130_fd_sc_hd__mux2i_4 _1077_ (.A0(_0748_),
    .A1(_0749_),
    .S(_0751_),
    .Y(_0752_));
 sky130_fd_sc_hd__clkinv_4 _1078_ (.A(_0752_),
    .Y(_0753_));
 sky130_fd_sc_hd__buf_4 _1079_ (.A(_0753_),
    .X(_0754_));
 sky130_fd_sc_hd__buf_4 _1080_ (.A(_0754_),
    .X(\compressed_decoder_i.instr_i[1] ));
 sky130_fd_sc_hd__mux2_2 _1081_ (.A0(net165),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[16] ),
    .S(_0746_),
    .X(_0755_));
 sky130_fd_sc_hd__mux2_1 _1082_ (.A0(net158),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[0] ),
    .S(_0746_),
    .X(_0756_));
 sky130_fd_sc_hd__mux2i_4 _1083_ (.A0(_0755_),
    .A1(_0756_),
    .S(_0751_),
    .Y(_0757_));
 sky130_fd_sc_hd__clkinv_8 _1084_ (.A(_0757_),
    .Y(_0758_));
 sky130_fd_sc_hd__buf_4 _1085_ (.A(_0758_),
    .X(\compressed_decoder_i.instr_i[0] ));
 sky130_fd_sc_hd__or2_1 _1086_ (.A(\gen_prefetch_buffer.prefetch_buffer_i.rdata_pmp_err_q[0] ),
    .B(net155),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_d[2] ));
 sky130_fd_sc_hd__buf_6 _1087_ (.A(_0751_),
    .X(_0759_));
 sky130_fd_sc_hd__nor2b_1 _1088_ (.A(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[0] ),
    .B_N(_0746_),
    .Y(_0760_));
 sky130_fd_sc_hd__nor3_1 _1089_ (.A(_0746_),
    .B(\gen_prefetch_buffer.prefetch_buffer_i.rdata_pmp_err_q[0] ),
    .C(net155),
    .Y(_0761_));
 sky130_fd_sc_hd__nand3_1 _1090_ (.A(_0747_),
    .B(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[16] ),
    .C(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[17] ),
    .Y(_0762_));
 sky130_fd_sc_hd__nand3b_1 _1091_ (.A_N(_0746_),
    .B(net165),
    .C(net166),
    .Y(_0763_));
 sky130_fd_sc_hd__o211ai_4 _1092_ (.A1(_0760_),
    .A2(_0761_),
    .B1(_0762_),
    .C1(_0763_),
    .Y(_0764_));
 sky130_fd_sc_hd__nand2_1 _1093_ (.A(net158),
    .B(net169),
    .Y(_0765_));
 sky130_fd_sc_hd__or2_1 _1094_ (.A(_0760_),
    .B(_0761_),
    .X(_0766_));
 sky130_fd_sc_hd__nand3_1 _1095_ (.A(_0747_),
    .B(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[0] ),
    .C(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[1] ),
    .Y(_0767_));
 sky130_fd_sc_hd__o2111ai_4 _1096_ (.A1(_0747_),
    .A2(_0765_),
    .B1(_0766_),
    .C1(_0751_),
    .D1(_0767_),
    .Y(_0768_));
 sky130_fd_sc_hd__o21ai_2 _1097_ (.A1(_0759_),
    .A2(_0764_),
    .B1(_0768_),
    .Y(_1060_));
 sky130_fd_sc_hd__inv_1 _1098_ (.A(_1060_),
    .Y(_1057_));
 sky130_fd_sc_hd__buf_2 _1099_ (.A(\gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .X(_0769_));
 sky130_fd_sc_hd__clkbuf_8 _1100_ (.A(net195),
    .X(_0770_));
 sky130_fd_sc_hd__buf_8 _1101_ (.A(_0770_),
    .X(_0771_));
 sky130_fd_sc_hd__buf_6 _1102_ (.A(pc_set_spec_i),
    .X(_0772_));
 sky130_fd_sc_hd__inv_2 _1103_ (.A(_0772_),
    .Y(_0773_));
 sky130_fd_sc_hd__buf_6 _1104_ (.A(net192),
    .X(_0774_));
 sky130_fd_sc_hd__nor2_4 _1105_ (.A(_0770_),
    .B(_0774_),
    .Y(_0775_));
 sky130_fd_sc_hd__buf_6 _1106_ (.A(\gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .X(_0776_));
 sky130_fd_sc_hd__o211ai_1 _1107_ (.A1(\gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ),
    .A2(\gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .B1(_0775_),
    .C1(_0776_),
    .Y(_0777_));
 sky130_fd_sc_hd__inv_1 _1108_ (.A(\gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1] ),
    .Y(_0778_));
 sky130_fd_sc_hd__o2111ai_1 _1109_ (.A1(_0771_),
    .A2(_0773_),
    .B1(net196),
    .C1(_0777_),
    .D1(_0778_),
    .Y(_0779_));
 sky130_fd_sc_hd__nand2b_1 _1110_ (.A_N(_0769_),
    .B(_0779_),
    .Y(_0780_));
 sky130_fd_sc_hd__buf_2 _1111_ (.A(_0780_),
    .X(net315));
 sky130_fd_sc_hd__inv_6 _1112_ (.A(net195),
    .Y(_0781_));
 sky130_fd_sc_hd__buf_8 _1113_ (.A(_0781_),
    .X(_0782_));
 sky130_fd_sc_hd__clkinv_2 _1114_ (.A(net192),
    .Y(_0783_));
 sky130_fd_sc_hd__buf_6 _1115_ (.A(_0783_),
    .X(_0784_));
 sky130_fd_sc_hd__nand2_8 _1116_ (.A(_0782_),
    .B(_0784_),
    .Y(_0785_));
 sky130_fd_sc_hd__o21a_1 _1117_ (.A1(\gen_prefetch_buffer.prefetch_buffer_i.discard_req_q ),
    .A2(_0785_),
    .B1(_0769_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.discard_req_d ));
 sky130_fd_sc_hd__mux2_2 _1118_ (.A0(net179),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[29] ),
    .S(_0745_),
    .X(_0786_));
 sky130_fd_sc_hd__mux2_1 _1119_ (.A0(net162),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[13] ),
    .S(_0745_),
    .X(_0787_));
 sky130_fd_sc_hd__mux2i_4 _1120_ (.A0(_0786_),
    .A1(_0787_),
    .S(_0750_),
    .Y(_0788_));
 sky130_fd_sc_hd__inv_1 _1121_ (.A(_0788_),
    .Y(_0789_));
 sky130_fd_sc_hd__buf_6 _1122_ (.A(_0789_),
    .X(_0790_));
 sky130_fd_sc_hd__buf_4 _1123_ (.A(_0790_),
    .X(_0791_));
 sky130_fd_sc_hd__buf_4 _1124_ (.A(_0791_),
    .X(\compressed_decoder_i.instr_i[13] ));
 sky130_fd_sc_hd__mux2_2 _1125_ (.A0(net181),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[30] ),
    .S(_0745_),
    .X(_0792_));
 sky130_fd_sc_hd__buf_6 _1126_ (.A(_0745_),
    .X(_0793_));
 sky130_fd_sc_hd__mux2_1 _1127_ (.A0(net163),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[14] ),
    .S(_0793_),
    .X(_0794_));
 sky130_fd_sc_hd__mux2i_4 _1128_ (.A0(_0792_),
    .A1(_0794_),
    .S(_0750_),
    .Y(_0795_));
 sky130_fd_sc_hd__inv_1 _1129_ (.A(_0795_),
    .Y(_0796_));
 sky130_fd_sc_hd__buf_6 _1130_ (.A(_0796_),
    .X(_0797_));
 sky130_fd_sc_hd__buf_6 _1131_ (.A(_0797_),
    .X(_0798_));
 sky130_fd_sc_hd__buf_4 _1132_ (.A(_0798_),
    .X(\compressed_decoder_i.instr_i[14] ));
 sky130_fd_sc_hd__buf_6 _1133_ (.A(net358),
    .X(_0799_));
 sky130_fd_sc_hd__mux4_4 _1134_ (.A0(net160),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[11] ),
    .A2(net177),
    .A3(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[27] ),
    .S0(_0793_),
    .S1(_0799_),
    .X(_0800_));
 sky130_fd_sc_hd__buf_6 _1135_ (.A(_0800_),
    .X(\compressed_decoder_i.instr_i[11] ));
 sky130_fd_sc_hd__mux4_4 _1136_ (.A0(net159),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[10] ),
    .A2(net176),
    .A3(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[26] ),
    .S0(_0745_),
    .S1(_0799_),
    .X(_0801_));
 sky130_fd_sc_hd__buf_4 _1137_ (.A(_0801_),
    .X(\compressed_decoder_i.instr_i[10] ));
 sky130_fd_sc_hd__mux4_4 _1138_ (.A0(net185),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[5] ),
    .A2(net171),
    .A3(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[21] ),
    .S0(_0793_),
    .S1(_0799_),
    .X(_0802_));
 sky130_fd_sc_hd__buf_4 _1139_ (.A(_0802_),
    .X(\compressed_decoder_i.instr_i[5] ));
 sky130_fd_sc_hd__mux4_4 _1140_ (.A0(net186),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[6] ),
    .A2(net172),
    .A3(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[22] ),
    .S0(_0793_),
    .S1(_0799_),
    .X(_0803_));
 sky130_fd_sc_hd__buf_4 _1141_ (.A(_0803_),
    .X(\compressed_decoder_i.instr_i[6] ));
 sky130_fd_sc_hd__mux2_2 _1142_ (.A0(net178),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[28] ),
    .S(_0793_),
    .X(_0804_));
 sky130_fd_sc_hd__mux2_1 _1143_ (.A0(net161),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[12] ),
    .S(_0793_),
    .X(_0805_));
 sky130_fd_sc_hd__mux2i_4 _1144_ (.A0(_0804_),
    .A1(_0805_),
    .S(_0750_),
    .Y(_0806_));
 sky130_fd_sc_hd__clkinv_2 _1145_ (.A(_0806_),
    .Y(_0807_));
 sky130_fd_sc_hd__buf_4 _1146_ (.A(_0807_),
    .X(_0808_));
 sky130_fd_sc_hd__buf_4 _1147_ (.A(_0808_),
    .X(\compressed_decoder_i.instr_i[12] ));
 sky130_fd_sc_hd__mux2i_4 _1148_ (.A0(net167),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[18] ),
    .S(_0747_),
    .Y(_0809_));
 sky130_fd_sc_hd__mux2i_2 _1149_ (.A0(net180),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[2] ),
    .S(_0747_),
    .Y(_0810_));
 sky130_fd_sc_hd__mux2i_4 _1150_ (.A0(_0809_),
    .A1(_0810_),
    .S(_0751_),
    .Y(_0811_));
 sky130_fd_sc_hd__buf_4 _1151_ (.A(_0811_),
    .X(\compressed_decoder_i.instr_i[2] ));
 sky130_fd_sc_hd__mux4_4 _1152_ (.A0(net183),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[3] ),
    .A2(net168),
    .A3(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[19] ),
    .S0(_0746_),
    .S1(_0799_),
    .X(\compressed_decoder_i.instr_i[3] ));
 sky130_fd_sc_hd__mux4_1 _1153_ (.A0(net184),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[4] ),
    .A2(net170),
    .A3(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[20] ),
    .S0(_0746_),
    .S1(_0799_),
    .X(_0812_));
 sky130_fd_sc_hd__buf_6 _1154_ (.A(_0812_),
    .X(\compressed_decoder_i.instr_i[4] ));
 sky130_fd_sc_hd__mux4_4 _1155_ (.A0(net187),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[7] ),
    .A2(net173),
    .A3(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[23] ),
    .S0(_0793_),
    .S1(_0799_),
    .X(_0813_));
 sky130_fd_sc_hd__buf_4 _1156_ (.A(_0813_),
    .X(\compressed_decoder_i.instr_i[7] ));
 sky130_fd_sc_hd__mux2_2 _1157_ (.A0(net174),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[24] ),
    .S(_0746_),
    .X(_0814_));
 sky130_fd_sc_hd__mux2_1 _1158_ (.A0(net188),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[8] ),
    .S(_0746_),
    .X(_0815_));
 sky130_fd_sc_hd__mux2i_4 _1159_ (.A0(_0814_),
    .A1(_0815_),
    .S(_0750_),
    .Y(_0816_));
 sky130_fd_sc_hd__clkinv_4 _1160_ (.A(_0816_),
    .Y(\compressed_decoder_i.instr_i[8] ));
 sky130_fd_sc_hd__mux2_2 _1161_ (.A0(net175),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[25] ),
    .S(_0745_),
    .X(_0817_));
 sky130_fd_sc_hd__mux2i_1 _1162_ (.A0(net189),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[9] ),
    .S(_0793_),
    .Y(_0818_));
 sky130_fd_sc_hd__nor2_1 _1163_ (.A(_0799_),
    .B(_0818_),
    .Y(_0819_));
 sky130_fd_sc_hd__a21oi_4 _1164_ (.A1(_0799_),
    .A2(_0817_),
    .B1(_0819_),
    .Y(_0820_));
 sky130_fd_sc_hd__clkinv_4 _1165_ (.A(_0820_),
    .Y(\compressed_decoder_i.instr_i[9] ));
 sky130_fd_sc_hd__buf_8 _1166_ (.A(_0776_),
    .X(_0821_));
 sky130_fd_sc_hd__mux2i_1 _1167_ (.A0(net183),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[35] ),
    .S(_0821_),
    .Y(_0822_));
 sky130_fd_sc_hd__inv_1 _1168_ (.A(_0822_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[3] ));
 sky130_fd_sc_hd__mux2_1 _1169_ (.A0(net184),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[36] ),
    .S(_0776_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[4] ));
 sky130_fd_sc_hd__mux2_1 _1170_ (.A0(net185),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[37] ),
    .S(_0821_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[5] ));
 sky130_fd_sc_hd__mux2i_1 _1171_ (.A0(net186),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[38] ),
    .S(_0776_),
    .Y(_0823_));
 sky130_fd_sc_hd__inv_1 _1172_ (.A(_0823_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[6] ));
 sky130_fd_sc_hd__mux2i_4 _1173_ (.A0(net187),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[39] ),
    .S(_0821_),
    .Y(_0824_));
 sky130_fd_sc_hd__inv_1 _1174_ (.A(_0824_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[7] ));
 sky130_fd_sc_hd__mux2_1 _1175_ (.A0(net188),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[40] ),
    .S(_0776_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[8] ));
 sky130_fd_sc_hd__mux2i_2 _1176_ (.A0(net189),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[41] ),
    .S(_0821_),
    .Y(_0825_));
 sky130_fd_sc_hd__inv_1 _1177_ (.A(_0825_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[9] ));
 sky130_fd_sc_hd__mux2i_1 _1178_ (.A0(net159),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[42] ),
    .S(_0776_),
    .Y(_0826_));
 sky130_fd_sc_hd__inv_1 _1179_ (.A(_0826_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[10] ));
 sky130_fd_sc_hd__mux2_1 _1180_ (.A0(net160),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[43] ),
    .S(_0776_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[11] ));
 sky130_fd_sc_hd__mux2i_2 _1181_ (.A0(net161),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[44] ),
    .S(_0821_),
    .Y(_0827_));
 sky130_fd_sc_hd__inv_1 _1182_ (.A(_0827_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[12] ));
 sky130_fd_sc_hd__mux2i_2 _1183_ (.A0(net162),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[45] ),
    .S(_0821_),
    .Y(_0828_));
 sky130_fd_sc_hd__inv_1 _1184_ (.A(_0828_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[13] ));
 sky130_fd_sc_hd__mux2_1 _1185_ (.A0(net163),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[46] ),
    .S(_0776_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[14] ));
 sky130_fd_sc_hd__mux2_1 _1186_ (.A0(net164),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[47] ),
    .S(_0821_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[15] ));
 sky130_fd_sc_hd__mux2_2 _1187_ (.A0(net182),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[31] ),
    .S(_0793_),
    .X(_0829_));
 sky130_fd_sc_hd__mux2_1 _1188_ (.A0(net164),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[15] ),
    .S(_0793_),
    .X(_0830_));
 sky130_fd_sc_hd__mux2i_4 _1189_ (.A0(_0829_),
    .A1(_0830_),
    .S(_0750_),
    .Y(_0831_));
 sky130_fd_sc_hd__inv_2 _1190_ (.A(_0831_),
    .Y(_0832_));
 sky130_fd_sc_hd__buf_6 _1191_ (.A(_0832_),
    .X(_0833_));
 sky130_fd_sc_hd__buf_4 _1192_ (.A(_0833_),
    .X(\compressed_decoder_i.instr_i[15] ));
 sky130_fd_sc_hd__buf_4 _1193_ (.A(_0774_),
    .X(_0834_));
 sky130_fd_sc_hd__buf_6 _1194_ (.A(_0834_),
    .X(_0835_));
 sky130_fd_sc_hd__buf_8 _1195_ (.A(_0799_),
    .X(_0836_));
 sky130_fd_sc_hd__and2_1 _1196_ (.A(_0836_),
    .B(_0764_),
    .X(_0837_));
 sky130_fd_sc_hd__o21ai_4 _1197_ (.A1(\gen_prefetch_buffer.prefetch_buffer_i.rdata_pmp_err_q[0] ),
    .A2(net190),
    .B1(\gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ),
    .Y(_0838_));
 sky130_fd_sc_hd__inv_1 _1198_ (.A(_0747_),
    .Y(_0839_));
 sky130_fd_sc_hd__o21ai_2 _1199_ (.A1(\gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0] ),
    .A2(_0838_),
    .B1(_0839_),
    .Y(_0840_));
 sky130_fd_sc_hd__clkinv_2 _1200_ (.A(\gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .Y(_0841_));
 sky130_fd_sc_hd__o31a_1 _1201_ (.A1(_0839_),
    .A2(\gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0] ),
    .A3(_0838_),
    .B1(_0841_),
    .X(_0842_));
 sky130_fd_sc_hd__nand3_2 _1202_ (.A(_0836_),
    .B(_0764_),
    .C(_0842_),
    .Y(_0843_));
 sky130_fd_sc_hd__o211ai_4 _1203_ (.A1(_0837_),
    .A2(_0840_),
    .B1(_0843_),
    .C1(net154),
    .Y(_0844_));
 sky130_fd_sc_hd__nor2_8 _1204_ (.A(_0835_),
    .B(_0844_),
    .Y(if_id_pipe_reg_we));
 sky130_fd_sc_hd__clkbuf_8 _1205_ (.A(\gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .X(_0845_));
 sky130_fd_sc_hd__buf_4 _1206_ (.A(_0845_),
    .X(_0846_));
 sky130_fd_sc_hd__nor4_4 _1207_ (.A(_0841_),
    .B(_0846_),
    .C(\gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0] ),
    .D(_0838_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[2] ));
 sky130_fd_sc_hd__buf_4 _1208_ (.A(net193),
    .X(_0847_));
 sky130_fd_sc_hd__clkinv_2 _1209_ (.A(_0847_),
    .Y(_0848_));
 sky130_fd_sc_hd__buf_4 _1210_ (.A(net194),
    .X(_0849_));
 sky130_fd_sc_hd__buf_4 _1211_ (.A(pc_mux_i[1]),
    .X(_0850_));
 sky130_fd_sc_hd__buf_8 _1212_ (.A(_0850_),
    .X(_0851_));
 sky130_fd_sc_hd__and3b_1 _1213_ (.A_N(_0849_),
    .B(_0851_),
    .C(net152),
    .X(_0852_));
 sky130_fd_sc_hd__buf_4 _1214_ (.A(net153),
    .X(_0853_));
 sky130_fd_sc_hd__or2_0 _1215_ (.A(_0853_),
    .B(net148),
    .X(_0854_));
 sky130_fd_sc_hd__nor3b_4 _1216_ (.A(_0851_),
    .B(_0847_),
    .C_N(_0849_),
    .Y(_0855_));
 sky130_fd_sc_hd__a32oi_4 _1217_ (.A1(_0848_),
    .A2(_0852_),
    .A3(_0854_),
    .B1(_0855_),
    .B2(net85),
    .Y(_0856_));
 sky130_fd_sc_hd__buf_6 _1218_ (.A(_0850_),
    .X(_0857_));
 sky130_fd_sc_hd__mux2i_2 _1219_ (.A0(net54),
    .A1(net116),
    .S(_0857_),
    .Y(_0858_));
 sky130_fd_sc_hd__nand2b_1 _1220_ (.A_N(net194),
    .B(net193),
    .Y(_0859_));
 sky130_fd_sc_hd__buf_8 _1221_ (.A(_0859_),
    .X(_0860_));
 sky130_fd_sc_hd__o21a_1 _1222_ (.A1(_0858_),
    .A2(_0860_),
    .B1(net195),
    .X(_0861_));
 sky130_fd_sc_hd__nor2b_1 _1223_ (.A(net192),
    .B_N(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[3] ),
    .Y(_0862_));
 sky130_fd_sc_hd__nor2_1 _1224_ (.A(_0770_),
    .B(_0862_),
    .Y(_0863_));
 sky130_fd_sc_hd__a21oi_2 _1225_ (.A1(_0856_),
    .A2(_0861_),
    .B1(_0863_),
    .Y(_1067_));
 sky130_fd_sc_hd__or2_4 _1226_ (.A(_0769_),
    .B(_0779_),
    .X(_0864_));
 sky130_fd_sc_hd__inv_1 _1227_ (.A(_0864_),
    .Y(_1064_));
 sky130_fd_sc_hd__clkbuf_4 _1228_ (.A(_0848_),
    .X(_0865_));
 sky130_fd_sc_hd__inv_1 _1229_ (.A(_0853_),
    .Y(_0866_));
 sky130_fd_sc_hd__and3_2 _1230_ (.A(_0865_),
    .B(_0866_),
    .C(_0852_),
    .X(_0867_));
 sky130_fd_sc_hd__buf_6 _1231_ (.A(_0860_),
    .X(_0868_));
 sky130_fd_sc_hd__buf_6 _1232_ (.A(_0857_),
    .X(_0869_));
 sky130_fd_sc_hd__buf_4 _1233_ (.A(_0869_),
    .X(_0870_));
 sky130_fd_sc_hd__mux2i_1 _1234_ (.A0(net51),
    .A1(net113),
    .S(_0870_),
    .Y(_0871_));
 sky130_fd_sc_hd__nor2_1 _1235_ (.A(_0868_),
    .B(_0871_),
    .Y(_0872_));
 sky130_fd_sc_hd__a221oi_4 _1236_ (.A1(net82),
    .A2(_0855_),
    .B1(_0867_),
    .B2(net147),
    .C1(_0872_),
    .Y(_0873_));
 sky130_fd_sc_hd__nand2_1 _1237_ (.A(_0784_),
    .B(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[2] ),
    .Y(_0874_));
 sky130_fd_sc_hd__buf_6 _1238_ (.A(_0782_),
    .X(_0875_));
 sky130_fd_sc_hd__mux2i_1 _1239_ (.A0(_0873_),
    .A1(_0874_),
    .S(_0875_),
    .Y(_1065_));
 sky130_fd_sc_hd__buf_4 _1240_ (.A(_0821_),
    .X(_0876_));
 sky130_fd_sc_hd__buf_4 _1241_ (.A(_0747_),
    .X(_0877_));
 sky130_fd_sc_hd__and3_1 _1242_ (.A(_0877_),
    .B(_0841_),
    .C(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_d[2] ),
    .X(_0878_));
 sky130_fd_sc_hd__a21oi_1 _1243_ (.A1(_0876_),
    .A2(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1] ),
    .B1(_0878_),
    .Y(_0879_));
 sky130_fd_sc_hd__nor3_1 _1244_ (.A(_0759_),
    .B(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[0] ),
    .C(_0879_),
    .Y(_0000_));
 sky130_fd_sc_hd__buf_4 _1245_ (.A(_0782_),
    .X(_0880_));
 sky130_fd_sc_hd__clkbuf_8 _1246_ (.A(_0880_),
    .X(_0881_));
 sky130_fd_sc_hd__buf_4 _1247_ (.A(net194),
    .X(_0882_));
 sky130_fd_sc_hd__buf_4 _1248_ (.A(_0882_),
    .X(_0883_));
 sky130_fd_sc_hd__buf_4 _1249_ (.A(_0883_),
    .X(_0884_));
 sky130_fd_sc_hd__or2_2 _1250_ (.A(_0851_),
    .B(_0847_),
    .X(_0885_));
 sky130_fd_sc_hd__nor3_2 _1251_ (.A(_0881_),
    .B(_0884_),
    .C(_0885_),
    .Y(net198));
 sky130_fd_sc_hd__a21boi_0 _1252_ (.A1(_0762_),
    .A2(_0763_),
    .B1_N(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_d[2] ),
    .Y(_0886_));
 sky130_fd_sc_hd__buf_6 _1253_ (.A(_0836_),
    .X(_0887_));
 sky130_fd_sc_hd__o21ai_0 _1254_ (.A1(_0876_),
    .A2(_0886_),
    .B1(_0887_),
    .Y(_0888_));
 sky130_fd_sc_hd__a2111oi_0 _1255_ (.A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1] ),
    .A2(_0764_),
    .B1(_0759_),
    .C1(_0841_),
    .D1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[0] ),
    .Y(_0889_));
 sky130_fd_sc_hd__a21oi_1 _1256_ (.A1(_0766_),
    .A2(_0888_),
    .B1(_0889_),
    .Y(fetch_err));
 sky130_fd_sc_hd__a21oi_1 _1257_ (.A1(\gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1] ),
    .A2(_0785_),
    .B1(\gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[1] ),
    .Y(_0890_));
 sky130_fd_sc_hd__or2_0 _1258_ (.A(net157),
    .B(net156),
    .X(_0891_));
 sky130_fd_sc_hd__buf_2 _1259_ (.A(_0891_),
    .X(_0892_));
 sky130_fd_sc_hd__clkbuf_2 _1260_ (.A(\gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ),
    .X(_0893_));
 sky130_fd_sc_hd__o21a_1 _1261_ (.A1(\gen_prefetch_buffer.prefetch_buffer_i.rdata_pmp_err_q[0] ),
    .A2(net190),
    .B1(_0893_),
    .X(_0894_));
 sky130_fd_sc_hd__a21oi_1 _1262_ (.A1(_0893_),
    .A2(_0785_),
    .B1(\gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0] ),
    .Y(_0895_));
 sky130_fd_sc_hd__nor2_1 _1263_ (.A(_0894_),
    .B(_0895_),
    .Y(_0896_));
 sky130_fd_sc_hd__a21oi_1 _1264_ (.A1(\gen_prefetch_buffer.prefetch_buffer_i.discard_req_d ),
    .A2(_0892_),
    .B1(_0896_),
    .Y(_0897_));
 sky130_fd_sc_hd__o21ai_0 _1265_ (.A1(_0838_),
    .A2(_0890_),
    .B1(_0897_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[0] ));
 sky130_fd_sc_hd__nand3_1 _1266_ (.A(_0893_),
    .B(\gen_prefetch_buffer.prefetch_buffer_i.discard_req_d ),
    .C(_0892_),
    .Y(_0898_));
 sky130_fd_sc_hd__a21oi_1 _1267_ (.A1(_0890_),
    .A2(_0898_),
    .B1(_0894_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[1] ));
 sky130_fd_sc_hd__buf_4 _1268_ (.A(_0771_),
    .X(_0899_));
 sky130_fd_sc_hd__buf_4 _1269_ (.A(_0849_),
    .X(_0900_));
 sky130_fd_sc_hd__nor2_8 _1270_ (.A(_0851_),
    .B(_0847_),
    .Y(_0901_));
 sky130_fd_sc_hd__buf_4 _1271_ (.A(net193),
    .X(_0902_));
 sky130_fd_sc_hd__nor3b_1 _1272_ (.A(_0902_),
    .B(_0853_),
    .C_N(net123),
    .Y(_0903_));
 sky130_fd_sc_hd__or3b_1 _1273_ (.A(_0850_),
    .B(net193),
    .C_N(net194),
    .X(_0904_));
 sky130_fd_sc_hd__o32a_2 _1274_ (.A1(_0900_),
    .A2(_0901_),
    .A3(_0903_),
    .B1(_0904_),
    .B2(net61),
    .X(_0905_));
 sky130_fd_sc_hd__buf_6 _1275_ (.A(_0857_),
    .X(_0906_));
 sky130_fd_sc_hd__mux2i_1 _1276_ (.A0(net30),
    .A1(net92),
    .S(_0906_),
    .Y(_0907_));
 sky130_fd_sc_hd__nor2_1 _1277_ (.A(_0868_),
    .B(_0907_),
    .Y(_0908_));
 sky130_fd_sc_hd__o21a_1 _1278_ (.A1(_0850_),
    .A2(net193),
    .B1(_0849_),
    .X(_0909_));
 sky130_fd_sc_hd__buf_6 _1279_ (.A(_0909_),
    .X(_0910_));
 sky130_fd_sc_hd__nor3_4 _1280_ (.A(_0849_),
    .B(_0851_),
    .C(_0902_),
    .Y(_0911_));
 sky130_fd_sc_hd__nor2_8 _1281_ (.A(_0910_),
    .B(_0911_),
    .Y(_0912_));
 sky130_fd_sc_hd__o22a_1 _1282_ (.A1(_0905_),
    .A2(_0908_),
    .B1(_0912_),
    .B2(net1),
    .X(_0913_));
 sky130_fd_sc_hd__buf_6 _1283_ (.A(_0770_),
    .X(_0914_));
 sky130_fd_sc_hd__nand2b_1 _1284_ (.A_N(_0774_),
    .B(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[10] ),
    .Y(_0915_));
 sky130_fd_sc_hd__nor2_1 _1285_ (.A(_0914_),
    .B(_0915_),
    .Y(_0916_));
 sky130_fd_sc_hd__a21oi_1 _1286_ (.A1(_0899_),
    .A2(_0913_),
    .B1(_0916_),
    .Y(_0917_));
 sky130_fd_sc_hd__or2_4 _1287_ (.A(_0849_),
    .B(_0847_),
    .X(_0918_));
 sky130_fd_sc_hd__buf_6 _1288_ (.A(_0851_),
    .X(_0919_));
 sky130_fd_sc_hd__clkinv_2 _1289_ (.A(_0919_),
    .Y(_0920_));
 sky130_fd_sc_hd__a21oi_1 _1290_ (.A1(_0866_),
    .A2(net145),
    .B1(_0920_),
    .Y(_0921_));
 sky130_fd_sc_hd__nor2b_1 _1291_ (.A(net121),
    .B_N(_0919_),
    .Y(_0922_));
 sky130_fd_sc_hd__inv_2 _1292_ (.A(_0882_),
    .Y(_0923_));
 sky130_fd_sc_hd__buf_4 _1293_ (.A(_0923_),
    .X(_0924_));
 sky130_fd_sc_hd__o21ai_1 _1294_ (.A1(_0865_),
    .A2(_0922_),
    .B1(_0924_),
    .Y(_0925_));
 sky130_fd_sc_hd__buf_4 _1295_ (.A(_0920_),
    .X(_0926_));
 sky130_fd_sc_hd__clkbuf_4 _1296_ (.A(_0847_),
    .X(_0927_));
 sky130_fd_sc_hd__o22ai_1 _1297_ (.A1(_0927_),
    .A2(net90),
    .B1(net59),
    .B2(_0883_),
    .Y(_0928_));
 sky130_fd_sc_hd__nand2_1 _1298_ (.A(_0926_),
    .B(_0928_),
    .Y(_0929_));
 sky130_fd_sc_hd__a2bb2oi_4 _1299_ (.A1_N(_0918_),
    .A2_N(_0921_),
    .B1(_0925_),
    .B2(_0929_),
    .Y(_0930_));
 sky130_fd_sc_hd__nor2_2 _1300_ (.A(net28),
    .B(_0912_),
    .Y(_0931_));
 sky130_fd_sc_hd__nor2b_4 _1301_ (.A(_0849_),
    .B_N(_0857_),
    .Y(_0932_));
 sky130_fd_sc_hd__nand2_2 _1302_ (.A(_0902_),
    .B(net120),
    .Y(_0933_));
 sky130_fd_sc_hd__nor4_2 _1303_ (.A(_0882_),
    .B(_0857_),
    .C(_0848_),
    .D(net58),
    .Y(_0934_));
 sky130_fd_sc_hd__nor2_2 _1304_ (.A(net89),
    .B(_0904_),
    .Y(_0935_));
 sky130_fd_sc_hd__a2111oi_4 _1305_ (.A1(_0932_),
    .A2(_0933_),
    .B1(_0934_),
    .C1(_0935_),
    .D1(_0781_),
    .Y(_0936_));
 sky130_fd_sc_hd__nor3b_4 _1306_ (.A(_0930_),
    .B(_0931_),
    .C_N(_0936_),
    .Y(_0937_));
 sky130_fd_sc_hd__and3_2 _1307_ (.A(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[7] ),
    .B(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[8] ),
    .C(_0775_),
    .X(_0938_));
 sky130_fd_sc_hd__mux2i_2 _1308_ (.A0(net55),
    .A1(net117),
    .S(_0919_),
    .Y(_0939_));
 sky130_fd_sc_hd__o2bb2ai_4 _1309_ (.A1_N(net86),
    .A2_N(_0855_),
    .B1(_0860_),
    .B2(_0939_),
    .Y(_0940_));
 sky130_fd_sc_hd__or4b_4 _1310_ (.A(net194),
    .B(net193),
    .C(net153),
    .D_N(_0850_),
    .X(_0941_));
 sky130_fd_sc_hd__nand2_1 _1311_ (.A(net152),
    .B(net149),
    .Y(_0942_));
 sky130_fd_sc_hd__o21ai_1 _1312_ (.A1(_0941_),
    .A2(_0942_),
    .B1(_0770_),
    .Y(_0943_));
 sky130_fd_sc_hd__nor2b_1 _1313_ (.A(net192),
    .B_N(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[4] ),
    .Y(_0944_));
 sky130_fd_sc_hd__or2_0 _1314_ (.A(net195),
    .B(_0944_),
    .X(_0945_));
 sky130_fd_sc_hd__o211ai_1 _1315_ (.A1(_0940_),
    .A2(_0943_),
    .B1(_0945_),
    .C1(_1068_),
    .Y(_0946_));
 sky130_fd_sc_hd__nor2b_1 _1316_ (.A(net192),
    .B_N(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[6] ),
    .Y(_0947_));
 sky130_fd_sc_hd__nand2_1 _1317_ (.A(net152),
    .B(net151),
    .Y(_0948_));
 sky130_fd_sc_hd__o21ai_2 _1318_ (.A1(_0941_),
    .A2(_0948_),
    .B1(_0770_),
    .Y(_0949_));
 sky130_fd_sc_hd__mux2i_1 _1319_ (.A0(net57),
    .A1(net119),
    .S(_0919_),
    .Y(_0950_));
 sky130_fd_sc_hd__o2bb2ai_2 _1320_ (.A1_N(net88),
    .A2_N(_0855_),
    .B1(_0860_),
    .B2(_0950_),
    .Y(_0951_));
 sky130_fd_sc_hd__o22ai_4 _1321_ (.A1(_0770_),
    .A2(_0947_),
    .B1(_0949_),
    .B2(_0951_),
    .Y(_0952_));
 sky130_fd_sc_hd__nor2b_1 _1322_ (.A(net192),
    .B_N(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[5] ),
    .Y(_0953_));
 sky130_fd_sc_hd__nand2_1 _1323_ (.A(net152),
    .B(net150),
    .Y(_0954_));
 sky130_fd_sc_hd__o21ai_2 _1324_ (.A1(_0941_),
    .A2(_0954_),
    .B1(net195),
    .Y(_0955_));
 sky130_fd_sc_hd__mux2i_1 _1325_ (.A0(net56),
    .A1(net118),
    .S(_0857_),
    .Y(_0956_));
 sky130_fd_sc_hd__o2bb2ai_2 _1326_ (.A1_N(net87),
    .A2_N(_0855_),
    .B1(_0860_),
    .B2(_0956_),
    .Y(_0957_));
 sky130_fd_sc_hd__o22ai_4 _1327_ (.A1(_0770_),
    .A2(_0953_),
    .B1(_0955_),
    .B2(_0957_),
    .Y(_0958_));
 sky130_fd_sc_hd__nor3_2 _1328_ (.A(_0946_),
    .B(_0952_),
    .C(_0958_),
    .Y(_0959_));
 sky130_fd_sc_hd__a21oi_1 _1329_ (.A1(_0866_),
    .A2(net146),
    .B1(_0926_),
    .Y(_0960_));
 sky130_fd_sc_hd__o22ai_1 _1330_ (.A1(_0927_),
    .A2(net91),
    .B1(net60),
    .B2(_0883_),
    .Y(_0961_));
 sky130_fd_sc_hd__nand2_1 _1331_ (.A(_0926_),
    .B(_0961_),
    .Y(_0962_));
 sky130_fd_sc_hd__nor2b_1 _1332_ (.A(net122),
    .B_N(_0906_),
    .Y(_0963_));
 sky130_fd_sc_hd__o21ai_1 _1333_ (.A1(_0865_),
    .A2(_0963_),
    .B1(_0924_),
    .Y(_0964_));
 sky130_fd_sc_hd__a2bb2oi_4 _1334_ (.A1_N(_0960_),
    .A2_N(_0918_),
    .B1(_0962_),
    .B2(_0964_),
    .Y(_0965_));
 sky130_fd_sc_hd__o21ai_2 _1335_ (.A1(net29),
    .A2(_0912_),
    .B1(_0771_),
    .Y(_0966_));
 sky130_fd_sc_hd__nand2_1 _1336_ (.A(_0784_),
    .B(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[9] ),
    .Y(_0967_));
 sky130_fd_sc_hd__o22ai_4 _1337_ (.A1(_0965_),
    .A2(_0966_),
    .B1(_0967_),
    .B2(_0771_),
    .Y(_0968_));
 sky130_fd_sc_hd__o211ai_4 _1338_ (.A1(_0937_),
    .A2(_0938_),
    .B1(_0959_),
    .C1(_0968_),
    .Y(_0969_));
 sky130_fd_sc_hd__buf_4 _1339_ (.A(_0969_),
    .X(_0970_));
 sky130_fd_sc_hd__xor2_1 _1340_ (.A(_0917_),
    .B(_0970_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[10] ));
 sky130_fd_sc_hd__nand2_1 _1341_ (.A(_0783_),
    .B(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[11] ),
    .Y(_0971_));
 sky130_fd_sc_hd__buf_4 _1342_ (.A(_0902_),
    .X(_0972_));
 sky130_fd_sc_hd__mux2i_1 _1343_ (.A0(net2),
    .A1(net31),
    .S(_0972_),
    .Y(_0973_));
 sky130_fd_sc_hd__nand3b_1 _1344_ (.A_N(_0972_),
    .B(net62),
    .C(_0900_),
    .Y(_0974_));
 sky130_fd_sc_hd__o21ai_2 _1345_ (.A1(_0883_),
    .A2(_0973_),
    .B1(_0974_),
    .Y(_0975_));
 sky130_fd_sc_hd__or3_1 _1346_ (.A(_0847_),
    .B(_0853_),
    .C(net124),
    .X(_0976_));
 sky130_fd_sc_hd__nand2b_1 _1347_ (.A_N(net93),
    .B(_0902_),
    .Y(_0977_));
 sky130_fd_sc_hd__a32o_1 _1348_ (.A1(_0932_),
    .A2(_0976_),
    .A3(_0977_),
    .B1(_0910_),
    .B2(net2),
    .X(_0978_));
 sky130_fd_sc_hd__a211oi_4 _1349_ (.A1(_0926_),
    .A2(_0975_),
    .B1(_0978_),
    .C1(_0781_),
    .Y(_0979_));
 sky130_fd_sc_hd__a21oi_1 _1350_ (.A1(_0880_),
    .A2(_0971_),
    .B1(_0979_),
    .Y(_0980_));
 sky130_fd_sc_hd__o211ai_2 _1351_ (.A1(_0940_),
    .A2(_0943_),
    .B1(_0945_),
    .C1(_1066_),
    .Y(_0981_));
 sky130_fd_sc_hd__nor4b_4 _1352_ (.A(_0952_),
    .B(_0958_),
    .C(_0981_),
    .D_N(_1067_),
    .Y(_0982_));
 sky130_fd_sc_hd__o211ai_4 _1353_ (.A1(_0937_),
    .A2(_0938_),
    .B1(_0982_),
    .C1(_0968_),
    .Y(_0983_));
 sky130_fd_sc_hd__buf_6 _1354_ (.A(_0983_),
    .X(_0984_));
 sky130_fd_sc_hd__nor2_1 _1355_ (.A(_0917_),
    .B(_0984_),
    .Y(_0985_));
 sky130_fd_sc_hd__xor2_1 _1356_ (.A(_0980_),
    .B(_0985_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[11] ));
 sky130_fd_sc_hd__nand2_1 _1357_ (.A(_0900_),
    .B(net3),
    .Y(_0986_));
 sky130_fd_sc_hd__mux2i_2 _1358_ (.A0(net32),
    .A1(net94),
    .S(_0906_),
    .Y(_0987_));
 sky130_fd_sc_hd__or4b_1 _1359_ (.A(_0882_),
    .B(_0857_),
    .C(_0902_),
    .D_N(net3),
    .X(_0988_));
 sky130_fd_sc_hd__o221ai_4 _1360_ (.A1(_0901_),
    .A2(_0986_),
    .B1(_0987_),
    .B2(_0860_),
    .C1(_0988_),
    .Y(_0989_));
 sky130_fd_sc_hd__nor2b_1 _1361_ (.A(net153),
    .B_N(_0851_),
    .Y(_0990_));
 sky130_fd_sc_hd__buf_4 _1362_ (.A(_0990_),
    .X(_0991_));
 sky130_fd_sc_hd__nor2b_1 _1363_ (.A(_0850_),
    .B_N(_0849_),
    .Y(_0992_));
 sky130_fd_sc_hd__buf_4 _1364_ (.A(_0992_),
    .X(_0993_));
 sky130_fd_sc_hd__a32o_1 _1365_ (.A1(_0924_),
    .A2(net125),
    .A3(_0991_),
    .B1(_0993_),
    .B2(net63),
    .X(_0994_));
 sky130_fd_sc_hd__buf_6 _1366_ (.A(_0972_),
    .X(_0995_));
 sky130_fd_sc_hd__nor2_2 _1367_ (.A(_0781_),
    .B(_0995_),
    .Y(_0996_));
 sky130_fd_sc_hd__nand2b_1 _1368_ (.A_N(_0774_),
    .B(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[12] ),
    .Y(_0997_));
 sky130_fd_sc_hd__nor2_1 _1369_ (.A(_0914_),
    .B(_0997_),
    .Y(_0998_));
 sky130_fd_sc_hd__a221oi_4 _1370_ (.A1(_0914_),
    .A2(_0989_),
    .B1(_0994_),
    .B2(_0996_),
    .C1(_0998_),
    .Y(_0999_));
 sky130_fd_sc_hd__o221ai_4 _1371_ (.A1(_0905_),
    .A2(_0908_),
    .B1(_0912_),
    .B2(net1),
    .C1(_0914_),
    .Y(_1000_));
 sky130_fd_sc_hd__inv_1 _1372_ (.A(_0916_),
    .Y(_1001_));
 sky130_fd_sc_hd__a221oi_4 _1373_ (.A1(_1000_),
    .A2(_1001_),
    .B1(_0971_),
    .B2(_0782_),
    .C1(_0979_),
    .Y(_1002_));
 sky130_fd_sc_hd__nor2b_1 _1374_ (.A(_0969_),
    .B_N(_1002_),
    .Y(_1003_));
 sky130_fd_sc_hd__xnor2_1 _1375_ (.A(_0999_),
    .B(_1003_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[12] ));
 sky130_fd_sc_hd__nand2_1 _1376_ (.A(_0883_),
    .B(net4),
    .Y(_1004_));
 sky130_fd_sc_hd__mux2i_2 _1377_ (.A0(net33),
    .A1(net95),
    .S(_0906_),
    .Y(_1005_));
 sky130_fd_sc_hd__or4b_1 _1378_ (.A(_0882_),
    .B(_0857_),
    .C(_0902_),
    .D_N(net4),
    .X(_1006_));
 sky130_fd_sc_hd__o221ai_4 _1379_ (.A1(_0901_),
    .A2(_1004_),
    .B1(_1005_),
    .B2(_0868_),
    .C1(_1006_),
    .Y(_1007_));
 sky130_fd_sc_hd__a32o_1 _1380_ (.A1(_0924_),
    .A2(net126),
    .A3(_0991_),
    .B1(_0993_),
    .B2(net64),
    .X(_1008_));
 sky130_fd_sc_hd__nand2b_1 _1381_ (.A_N(_0774_),
    .B(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[13] ),
    .Y(_1009_));
 sky130_fd_sc_hd__nor2_1 _1382_ (.A(_0914_),
    .B(_1009_),
    .Y(_1010_));
 sky130_fd_sc_hd__a221oi_4 _1383_ (.A1(_0771_),
    .A2(_1007_),
    .B1(_1008_),
    .B2(_0996_),
    .C1(_1010_),
    .Y(_1011_));
 sky130_fd_sc_hd__nor3b_1 _1384_ (.A(_0984_),
    .B(_0999_),
    .C_N(_1002_),
    .Y(_1012_));
 sky130_fd_sc_hd__xnor2_1 _1385_ (.A(_1011_),
    .B(_1012_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[13] ));
 sky130_fd_sc_hd__nand2b_1 _1386_ (.A_N(_0853_),
    .B(net127),
    .Y(_1013_));
 sky130_fd_sc_hd__a21oi_2 _1387_ (.A1(_0869_),
    .A2(_1013_),
    .B1(_0918_),
    .Y(_1014_));
 sky130_fd_sc_hd__mux2i_1 _1388_ (.A0(net34),
    .A1(net96),
    .S(_0906_),
    .Y(_1015_));
 sky130_fd_sc_hd__o2bb2ai_1 _1389_ (.A1_N(net65),
    .A2_N(_0855_),
    .B1(_0868_),
    .B2(_1015_),
    .Y(_1016_));
 sky130_fd_sc_hd__o32ai_4 _1390_ (.A1(_0910_),
    .A2(_1014_),
    .A3(_1016_),
    .B1(_0912_),
    .B2(net5),
    .Y(_1017_));
 sky130_fd_sc_hd__nand3_1 _1391_ (.A(_0782_),
    .B(_0784_),
    .C(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[14] ),
    .Y(_1018_));
 sky130_fd_sc_hd__o21ai_4 _1392_ (.A1(_0782_),
    .A2(_1017_),
    .B1(_1018_),
    .Y(_1019_));
 sky130_fd_sc_hd__nor2_2 _1393_ (.A(_0999_),
    .B(_1011_),
    .Y(_1020_));
 sky130_fd_sc_hd__nand2_1 _1394_ (.A(_1002_),
    .B(_1020_),
    .Y(_1021_));
 sky130_fd_sc_hd__nor2_1 _1395_ (.A(_0970_),
    .B(_1021_),
    .Y(_1022_));
 sky130_fd_sc_hd__xor2_1 _1396_ (.A(_1019_),
    .B(_1022_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[14] ));
 sky130_fd_sc_hd__nand3_4 _1397_ (.A(_1002_),
    .B(_1019_),
    .C(_1020_),
    .Y(_1023_));
 sky130_fd_sc_hd__nor2_1 _1398_ (.A(_0984_),
    .B(_1023_),
    .Y(_1024_));
 sky130_fd_sc_hd__nand3b_1 _1399_ (.A_N(_0857_),
    .B(net66),
    .C(_0882_),
    .Y(_1025_));
 sky130_fd_sc_hd__nand4bb_1 _1400_ (.A_N(net194),
    .B_N(net153),
    .C(net128),
    .D(_0850_),
    .Y(_1026_));
 sky130_fd_sc_hd__a21oi_2 _1401_ (.A1(_1025_),
    .A2(_1026_),
    .B1(_0927_),
    .Y(_1027_));
 sky130_fd_sc_hd__and3_1 _1402_ (.A(_0882_),
    .B(net11),
    .C(_0885_),
    .X(_1028_));
 sky130_fd_sc_hd__and3_1 _1403_ (.A(_0923_),
    .B(net11),
    .C(_0901_),
    .X(_1029_));
 sky130_fd_sc_hd__mux2i_1 _1404_ (.A0(net35),
    .A1(net97),
    .S(_0919_),
    .Y(_1030_));
 sky130_fd_sc_hd__nor2_1 _1405_ (.A(_0860_),
    .B(_1030_),
    .Y(_1031_));
 sky130_fd_sc_hd__o41ai_4 _1406_ (.A1(_1027_),
    .A2(_1028_),
    .A3(_1029_),
    .A4(_1031_),
    .B1(_0914_),
    .Y(_1032_));
 sky130_fd_sc_hd__buf_6 _1407_ (.A(_0775_),
    .X(_1033_));
 sky130_fd_sc_hd__nand2_1 _1408_ (.A(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[15] ),
    .B(_1033_),
    .Y(_1034_));
 sky130_fd_sc_hd__nand2_1 _1409_ (.A(_1032_),
    .B(_1034_),
    .Y(_1035_));
 sky130_fd_sc_hd__xor2_1 _1410_ (.A(_1024_),
    .B(_1035_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[15] ));
 sky130_fd_sc_hd__a21oi_1 _1411_ (.A1(_0865_),
    .A2(net12),
    .B1(_0869_),
    .Y(_1036_));
 sky130_fd_sc_hd__or3_1 _1412_ (.A(_0902_),
    .B(_0853_),
    .C(net129),
    .X(_1037_));
 sky130_fd_sc_hd__o221ai_1 _1413_ (.A1(_0848_),
    .A2(net98),
    .B1(_1037_),
    .B2(_0926_),
    .C1(_0924_),
    .Y(_1038_));
 sky130_fd_sc_hd__nor4bb_1 _1414_ (.A(_0882_),
    .B(_0919_),
    .C_N(_0972_),
    .D_N(net36),
    .Y(_1039_));
 sky130_fd_sc_hd__a31oi_1 _1415_ (.A1(_0865_),
    .A2(net67),
    .A3(_0993_),
    .B1(_1039_),
    .Y(_1040_));
 sky130_fd_sc_hd__nand2_1 _1416_ (.A(net12),
    .B(_0910_),
    .Y(_1041_));
 sky130_fd_sc_hd__o211a_2 _1417_ (.A1(_1036_),
    .A2(_1038_),
    .B1(_1040_),
    .C1(_1041_),
    .X(_1042_));
 sky130_fd_sc_hd__nor2_2 _1418_ (.A(_0880_),
    .B(_1042_),
    .Y(_1043_));
 sky130_fd_sc_hd__a21oi_1 _1419_ (.A1(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[16] ),
    .A2(_1033_),
    .B1(_1043_),
    .Y(_1044_));
 sky130_fd_sc_hd__nor3b_1 _1420_ (.A(_0970_),
    .B(_1023_),
    .C_N(_1035_),
    .Y(_1045_));
 sky130_fd_sc_hd__xnor2_1 _1421_ (.A(_1044_),
    .B(_1045_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[16] ));
 sky130_fd_sc_hd__nor2_1 _1422_ (.A(_1032_),
    .B(_1042_),
    .Y(_1046_));
 sky130_fd_sc_hd__a31oi_1 _1423_ (.A1(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[15] ),
    .A2(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[16] ),
    .A3(_1033_),
    .B1(_1046_),
    .Y(_1047_));
 sky130_fd_sc_hd__nor3_1 _1424_ (.A(_0984_),
    .B(_1023_),
    .C(_1047_),
    .Y(_1048_));
 sky130_fd_sc_hd__or2_0 _1425_ (.A(_0910_),
    .B(_0911_),
    .X(_1049_));
 sky130_fd_sc_hd__mux2_1 _1426_ (.A0(net37),
    .A1(net99),
    .S(_0919_),
    .X(_1050_));
 sky130_fd_sc_hd__nor2b_4 _1427_ (.A(_0900_),
    .B_N(_0972_),
    .Y(_1051_));
 sky130_fd_sc_hd__a32o_1 _1428_ (.A1(_0923_),
    .A2(net130),
    .A3(_0991_),
    .B1(_0993_),
    .B2(net68),
    .X(_1052_));
 sky130_fd_sc_hd__a222oi_1 _1429_ (.A1(net13),
    .A2(_1049_),
    .B1(_1050_),
    .B2(_1051_),
    .C1(_1052_),
    .C2(_0865_),
    .Y(_1053_));
 sky130_fd_sc_hd__nand2_1 _1430_ (.A(_0784_),
    .B(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[17] ),
    .Y(_1054_));
 sky130_fd_sc_hd__mux2i_1 _1431_ (.A0(net8),
    .A1(_1054_),
    .S(_0880_),
    .Y(_1055_));
 sky130_fd_sc_hd__xor2_1 _1432_ (.A(_1048_),
    .B(_1055_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[17] ));
 sky130_fd_sc_hd__nand4_1 _1433_ (.A(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[15] ),
    .B(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[16] ),
    .C(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[17] ),
    .D(_0775_),
    .Y(_0001_));
 sky130_fd_sc_hd__o31ai_4 _1434_ (.A1(_1032_),
    .A2(_1042_),
    .A3(net8),
    .B1(_0001_),
    .Y(_0002_));
 sky130_fd_sc_hd__nand4_2 _1435_ (.A(_1002_),
    .B(_1019_),
    .C(_1020_),
    .D(_0002_),
    .Y(_0003_));
 sky130_fd_sc_hd__nor2_1 _1436_ (.A(_0970_),
    .B(_0003_),
    .Y(_0004_));
 sky130_fd_sc_hd__inv_2 _1437_ (.A(net14),
    .Y(_0005_));
 sky130_fd_sc_hd__a32oi_4 _1438_ (.A1(_0924_),
    .A2(net131),
    .A3(_0991_),
    .B1(_0993_),
    .B2(net69),
    .Y(_0006_));
 sky130_fd_sc_hd__mux2_1 _1439_ (.A0(net38),
    .A1(net100),
    .S(_0906_),
    .X(_0007_));
 sky130_fd_sc_hd__nand2_1 _1440_ (.A(_1051_),
    .B(_0007_),
    .Y(_0008_));
 sky130_fd_sc_hd__o221ai_4 _1441_ (.A1(_0005_),
    .A2(_0912_),
    .B1(_0006_),
    .B2(_0995_),
    .C1(_0008_),
    .Y(_0009_));
 sky130_fd_sc_hd__nand2_1 _1442_ (.A(_0784_),
    .B(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[18] ),
    .Y(_0010_));
 sky130_fd_sc_hd__nor2_1 _1443_ (.A(_0899_),
    .B(_0010_),
    .Y(_0011_));
 sky130_fd_sc_hd__a21o_1 _1444_ (.A1(_0899_),
    .A2(_0009_),
    .B1(_0011_),
    .X(_0012_));
 sky130_fd_sc_hd__xor2_1 _1445_ (.A(_0004_),
    .B(_0012_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[18] ));
 sky130_fd_sc_hd__mux2i_2 _1446_ (.A0(net39),
    .A1(net101),
    .S(_0869_),
    .Y(_0013_));
 sky130_fd_sc_hd__a32oi_4 _1447_ (.A1(_0924_),
    .A2(net132),
    .A3(_0991_),
    .B1(_0993_),
    .B2(net70),
    .Y(_0014_));
 sky130_fd_sc_hd__o21ai_2 _1448_ (.A1(_0910_),
    .A2(_0911_),
    .B1(net15),
    .Y(_0015_));
 sky130_fd_sc_hd__o221ai_4 _1449_ (.A1(_0868_),
    .A2(_0013_),
    .B1(_0014_),
    .B2(_0995_),
    .C1(_0015_),
    .Y(_0016_));
 sky130_fd_sc_hd__buf_4 _1450_ (.A(_0899_),
    .X(_0017_));
 sky130_fd_sc_hd__a22oi_1 _1451_ (.A1(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[19] ),
    .A2(_1033_),
    .B1(_0016_),
    .B2(_0017_),
    .Y(_0018_));
 sky130_fd_sc_hd__nand2_1 _1452_ (.A(_0002_),
    .B(_0012_),
    .Y(_0019_));
 sky130_fd_sc_hd__nor3_1 _1453_ (.A(_0984_),
    .B(_1023_),
    .C(_0019_),
    .Y(_0020_));
 sky130_fd_sc_hd__xnor2_1 _1454_ (.A(_0018_),
    .B(_0020_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[19] ));
 sky130_fd_sc_hd__nand3b_1 _1455_ (.A_N(_0900_),
    .B(_0927_),
    .C(net41),
    .Y(_0021_));
 sky130_fd_sc_hd__nand3b_1 _1456_ (.A_N(_0927_),
    .B(net72),
    .C(_0883_),
    .Y(_0022_));
 sky130_fd_sc_hd__a21oi_1 _1457_ (.A1(_0021_),
    .A2(_0022_),
    .B1(_0869_),
    .Y(_0023_));
 sky130_fd_sc_hd__or3_1 _1458_ (.A(_0902_),
    .B(_0853_),
    .C(net133),
    .X(_0024_));
 sky130_fd_sc_hd__o211a_1 _1459_ (.A1(_0848_),
    .A2(net103),
    .B1(_0932_),
    .C1(_0024_),
    .X(_0025_));
 sky130_fd_sc_hd__a211o_2 _1460_ (.A1(net16),
    .A2(_1049_),
    .B1(_0023_),
    .C1(_0025_),
    .X(_0026_));
 sky130_fd_sc_hd__a22oi_1 _1461_ (.A1(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[20] ),
    .A2(_1033_),
    .B1(_0026_),
    .B2(_0017_),
    .Y(_0027_));
 sky130_fd_sc_hd__nor3b_1 _1462_ (.A(_0010_),
    .B(_0899_),
    .C_N(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[19] ),
    .Y(_0028_));
 sky130_fd_sc_hd__a31oi_1 _1463_ (.A1(_0017_),
    .A2(_0009_),
    .A3(_0016_),
    .B1(_0028_),
    .Y(_0029_));
 sky130_fd_sc_hd__nor3_1 _1464_ (.A(_0970_),
    .B(_0003_),
    .C(_0029_),
    .Y(_0030_));
 sky130_fd_sc_hd__xnor2_1 _1465_ (.A(_0027_),
    .B(_0030_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[20] ));
 sky130_fd_sc_hd__nor4b_4 _1466_ (.A(_0900_),
    .B(_0972_),
    .C(_0853_),
    .D_N(_0919_),
    .Y(_0031_));
 sky130_fd_sc_hd__mux2i_1 _1467_ (.A0(net42),
    .A1(net104),
    .S(_0869_),
    .Y(_0032_));
 sky130_fd_sc_hd__o2bb2ai_2 _1468_ (.A1_N(net134),
    .A2_N(_0031_),
    .B1(_0032_),
    .B2(_0868_),
    .Y(_0033_));
 sky130_fd_sc_hd__or4b_1 _1469_ (.A(_0900_),
    .B(_0906_),
    .C(_0972_),
    .D_N(net17),
    .X(_0034_));
 sky130_fd_sc_hd__or4bb_1 _1470_ (.A(_0906_),
    .B(_0972_),
    .C_N(net73),
    .D_N(_0900_),
    .X(_0035_));
 sky130_fd_sc_hd__o211ai_1 _1471_ (.A1(_0870_),
    .A2(_0995_),
    .B1(net17),
    .C1(_0884_),
    .Y(_0036_));
 sky130_fd_sc_hd__nand3_2 _1472_ (.A(_0034_),
    .B(_0035_),
    .C(_0036_),
    .Y(_0037_));
 sky130_fd_sc_hd__o21ai_4 _1473_ (.A1(_0033_),
    .A2(_0037_),
    .B1(_0771_),
    .Y(_0038_));
 sky130_fd_sc_hd__nand2_1 _1474_ (.A(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[21] ),
    .B(_1033_),
    .Y(_0039_));
 sky130_fd_sc_hd__nand2_1 _1475_ (.A(_0038_),
    .B(_0039_),
    .Y(_0040_));
 sky130_fd_sc_hd__and4_1 _1476_ (.A(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[18] ),
    .B(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[19] ),
    .C(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[20] ),
    .D(_0775_),
    .X(_0041_));
 sky130_fd_sc_hd__a41o_1 _1477_ (.A1(_0771_),
    .A2(_0009_),
    .A3(_0016_),
    .A4(_0026_),
    .B1(_0041_),
    .X(_0042_));
 sky130_fd_sc_hd__nor3b_1 _1478_ (.A(_0984_),
    .B(_0003_),
    .C_N(_0042_),
    .Y(_0043_));
 sky130_fd_sc_hd__xor2_1 _1479_ (.A(_0040_),
    .B(_0043_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[21] ));
 sky130_fd_sc_hd__buf_4 _1480_ (.A(_0017_),
    .X(_0044_));
 sky130_fd_sc_hd__nor2b_1 _1481_ (.A(_0774_),
    .B_N(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[22] ),
    .Y(_0045_));
 sky130_fd_sc_hd__mux2_1 _1482_ (.A0(net18),
    .A1(net74),
    .S(_0901_),
    .X(_0046_));
 sky130_fd_sc_hd__and3_1 _1483_ (.A(_0924_),
    .B(net18),
    .C(_0901_),
    .X(_0047_));
 sky130_fd_sc_hd__mux2i_1 _1484_ (.A0(net43),
    .A1(net105),
    .S(_0870_),
    .Y(_0048_));
 sky130_fd_sc_hd__o2bb2ai_1 _1485_ (.A1_N(net135),
    .A2_N(_0031_),
    .B1(_0048_),
    .B2(_0868_),
    .Y(_0049_));
 sky130_fd_sc_hd__a211oi_4 _1486_ (.A1(_0884_),
    .A2(_0046_),
    .B1(_0047_),
    .C1(_0049_),
    .Y(_0050_));
 sky130_fd_sc_hd__and2_2 _1487_ (.A(_0899_),
    .B(_0050_),
    .X(_0051_));
 sky130_fd_sc_hd__o21bai_1 _1488_ (.A1(_0044_),
    .A2(_0045_),
    .B1_N(_0051_),
    .Y(_0052_));
 sky130_fd_sc_hd__nand2_1 _1489_ (.A(_0040_),
    .B(_0042_),
    .Y(_0053_));
 sky130_fd_sc_hd__or3_1 _1490_ (.A(_0969_),
    .B(_0003_),
    .C(_0053_),
    .X(_0054_));
 sky130_fd_sc_hd__nand3_1 _1491_ (.A(_0782_),
    .B(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[21] ),
    .C(_0045_),
    .Y(_0055_));
 sky130_fd_sc_hd__a22oi_2 _1492_ (.A1(_0899_),
    .A2(_0050_),
    .B1(_0055_),
    .B2(_0038_),
    .Y(_0056_));
 sky130_fd_sc_hd__nand3_2 _1493_ (.A(_0002_),
    .B(_0042_),
    .C(_0056_),
    .Y(_0057_));
 sky130_fd_sc_hd__nor3_1 _1494_ (.A(_0970_),
    .B(_1023_),
    .C(_0057_),
    .Y(_0058_));
 sky130_fd_sc_hd__a21oi_1 _1495_ (.A1(_0052_),
    .A2(_0054_),
    .B1(_0058_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[22] ));
 sky130_fd_sc_hd__nand2b_1 _1496_ (.A_N(net153),
    .B(net136),
    .Y(_0059_));
 sky130_fd_sc_hd__a21oi_2 _1497_ (.A1(_0919_),
    .A2(_0059_),
    .B1(_0918_),
    .Y(_0060_));
 sky130_fd_sc_hd__mux2i_1 _1498_ (.A0(net44),
    .A1(net106),
    .S(_0857_),
    .Y(_0061_));
 sky130_fd_sc_hd__o2bb2ai_2 _1499_ (.A1_N(net75),
    .A2_N(_0855_),
    .B1(_0860_),
    .B2(_0061_),
    .Y(_0062_));
 sky130_fd_sc_hd__o21bai_2 _1500_ (.A1(_0910_),
    .A2(_0911_),
    .B1_N(net19),
    .Y(_0063_));
 sky130_fd_sc_hd__o311ai_4 _1501_ (.A1(_0910_),
    .A2(_0060_),
    .A3(_0062_),
    .B1(_0063_),
    .C1(_0914_),
    .Y(_0064_));
 sky130_fd_sc_hd__nand3_2 _1502_ (.A(_0782_),
    .B(_0783_),
    .C(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[23] ),
    .Y(_0065_));
 sky130_fd_sc_hd__nand2_1 _1503_ (.A(_0064_),
    .B(_0065_),
    .Y(_0066_));
 sky130_fd_sc_hd__nor3_1 _1504_ (.A(_0984_),
    .B(_1023_),
    .C(_0057_),
    .Y(_0067_));
 sky130_fd_sc_hd__xor2_1 _1505_ (.A(_0066_),
    .B(_0067_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[23] ));
 sky130_fd_sc_hd__nand2_1 _1506_ (.A(_0882_),
    .B(net20),
    .Y(_0068_));
 sky130_fd_sc_hd__mux2i_1 _1507_ (.A0(net45),
    .A1(net107),
    .S(_0851_),
    .Y(_0069_));
 sky130_fd_sc_hd__or4b_1 _1508_ (.A(net194),
    .B(_0850_),
    .C(net193),
    .D_N(net20),
    .X(_0070_));
 sky130_fd_sc_hd__o221a_2 _1509_ (.A1(_0901_),
    .A2(_0068_),
    .B1(_0069_),
    .B2(_0860_),
    .C1(_0070_),
    .X(_0071_));
 sky130_fd_sc_hd__a32oi_4 _1510_ (.A1(_0923_),
    .A2(net137),
    .A3(_0991_),
    .B1(_0993_),
    .B2(net76),
    .Y(_0072_));
 sky130_fd_sc_hd__nand2_1 _1511_ (.A(_0770_),
    .B(_0865_),
    .Y(_0073_));
 sky130_fd_sc_hd__nand3_1 _1512_ (.A(_0781_),
    .B(_0783_),
    .C(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[24] ),
    .Y(_0074_));
 sky130_fd_sc_hd__o221a_2 _1513_ (.A1(_0781_),
    .A2(_0071_),
    .B1(_0072_),
    .B2(_0073_),
    .C1(_0074_),
    .X(_0075_));
 sky130_fd_sc_hd__nand3_2 _1514_ (.A(_1002_),
    .B(_1020_),
    .C(_0002_),
    .Y(_0076_));
 sky130_fd_sc_hd__nand3_2 _1515_ (.A(_1019_),
    .B(_0042_),
    .C(_0056_),
    .Y(_0077_));
 sky130_fd_sc_hd__nor4b_1 _1516_ (.A(_0970_),
    .B(_0076_),
    .C(_0077_),
    .D_N(_0066_),
    .Y(_0078_));
 sky130_fd_sc_hd__xnor2_1 _1517_ (.A(_0075_),
    .B(_0078_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[24] ));
 sky130_fd_sc_hd__mux2_1 _1518_ (.A0(net21),
    .A1(net46),
    .S(_0847_),
    .X(_0079_));
 sky130_fd_sc_hd__nand2_1 _1519_ (.A(_0906_),
    .B(_0972_),
    .Y(_0080_));
 sky130_fd_sc_hd__o221ai_1 _1520_ (.A1(_0906_),
    .A2(_0079_),
    .B1(_0080_),
    .B2(net108),
    .C1(_0923_),
    .Y(_0081_));
 sky130_fd_sc_hd__or3_1 _1521_ (.A(_0851_),
    .B(_0847_),
    .C(net77),
    .X(_0082_));
 sky130_fd_sc_hd__nand2b_1 _1522_ (.A_N(net21),
    .B(_0902_),
    .Y(_0083_));
 sky130_fd_sc_hd__a31oi_1 _1523_ (.A1(_0883_),
    .A2(_0082_),
    .A3(_0083_),
    .B1(_0781_),
    .Y(_0084_));
 sky130_fd_sc_hd__a21oi_2 _1524_ (.A1(_0783_),
    .A2(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[25] ),
    .B1(_0770_),
    .Y(_0085_));
 sky130_fd_sc_hd__nand2b_1 _1525_ (.A_N(net21),
    .B(_0882_),
    .Y(_0086_));
 sky130_fd_sc_hd__or4_1 _1526_ (.A(_0849_),
    .B(net193),
    .C(net153),
    .D(net138),
    .X(_0087_));
 sky130_fd_sc_hd__a211oi_1 _1527_ (.A1(_0086_),
    .A2(_0087_),
    .B1(_0781_),
    .C1(_0926_),
    .Y(_0088_));
 sky130_fd_sc_hd__a211o_2 _1528_ (.A1(_0081_),
    .A2(_0084_),
    .B1(_0085_),
    .C1(_0088_),
    .X(_0089_));
 sky130_fd_sc_hd__a21oi_1 _1529_ (.A1(_0064_),
    .A2(_0065_),
    .B1(_0075_),
    .Y(_0090_));
 sky130_fd_sc_hd__nor4b_1 _1530_ (.A(_0984_),
    .B(_0076_),
    .C(_0077_),
    .D_N(_0090_),
    .Y(_0091_));
 sky130_fd_sc_hd__xnor2_1 _1531_ (.A(_0089_),
    .B(_0091_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[25] ));
 sky130_fd_sc_hd__nand2_1 _1532_ (.A(_0900_),
    .B(net22),
    .Y(_0092_));
 sky130_fd_sc_hd__mux2i_2 _1533_ (.A0(net47),
    .A1(net109),
    .S(_0919_),
    .Y(_0093_));
 sky130_fd_sc_hd__or4b_1 _1534_ (.A(_0849_),
    .B(_0851_),
    .C(_0847_),
    .D_N(net22),
    .X(_0094_));
 sky130_fd_sc_hd__o221ai_4 _1535_ (.A1(_0901_),
    .A2(_0092_),
    .B1(_0093_),
    .B2(_0860_),
    .C1(_0094_),
    .Y(_0095_));
 sky130_fd_sc_hd__a32o_1 _1536_ (.A1(_0923_),
    .A2(net139),
    .A3(_0991_),
    .B1(_0993_),
    .B2(net78),
    .X(_0096_));
 sky130_fd_sc_hd__nand2b_1 _1537_ (.A_N(_0774_),
    .B(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[26] ),
    .Y(_0097_));
 sky130_fd_sc_hd__nor2_1 _1538_ (.A(_0914_),
    .B(_0097_),
    .Y(_0098_));
 sky130_fd_sc_hd__a221oi_4 _1539_ (.A1(_0914_),
    .A2(_0095_),
    .B1(_0096_),
    .B2(_0996_),
    .C1(_0098_),
    .Y(_0099_));
 sky130_fd_sc_hd__nor2b_1 _1540_ (.A(_0089_),
    .B_N(_0090_),
    .Y(_0100_));
 sky130_fd_sc_hd__nor4b_1 _1541_ (.A(_0970_),
    .B(_0076_),
    .C(_0077_),
    .D_N(_0100_),
    .Y(_0101_));
 sky130_fd_sc_hd__xnor2_1 _1542_ (.A(_0099_),
    .B(_0101_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[26] ));
 sky130_fd_sc_hd__a21oi_1 _1543_ (.A1(_0784_),
    .A2(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[27] ),
    .B1(_0771_),
    .Y(_0102_));
 sky130_fd_sc_hd__mux2i_1 _1544_ (.A0(net23),
    .A1(net48),
    .S(_0995_),
    .Y(_0103_));
 sky130_fd_sc_hd__nand3b_1 _1545_ (.A_N(_0995_),
    .B(net79),
    .C(_0883_),
    .Y(_0104_));
 sky130_fd_sc_hd__o21ai_2 _1546_ (.A1(_0884_),
    .A2(_0103_),
    .B1(_0104_),
    .Y(_0105_));
 sky130_fd_sc_hd__or3_1 _1547_ (.A(_0972_),
    .B(_0853_),
    .C(net140),
    .X(_0106_));
 sky130_fd_sc_hd__nand2b_1 _1548_ (.A_N(net110),
    .B(_0927_),
    .Y(_0107_));
 sky130_fd_sc_hd__a32o_1 _1549_ (.A1(_0932_),
    .A2(_0106_),
    .A3(_0107_),
    .B1(_0910_),
    .B2(net23),
    .X(_0108_));
 sky130_fd_sc_hd__a211oi_4 _1550_ (.A1(_0926_),
    .A2(_0105_),
    .B1(_0108_),
    .C1(_0782_),
    .Y(_0109_));
 sky130_fd_sc_hd__nor2_1 _1551_ (.A(_0102_),
    .B(_0109_),
    .Y(_0110_));
 sky130_fd_sc_hd__a2111oi_4 _1552_ (.A1(_0064_),
    .A2(_0065_),
    .B1(_0075_),
    .C1(_0089_),
    .D1(_0099_),
    .Y(_0111_));
 sky130_fd_sc_hd__nor4b_1 _1553_ (.A(_0983_),
    .B(_1023_),
    .C(_0057_),
    .D_N(_0111_),
    .Y(_0112_));
 sky130_fd_sc_hd__xor2_1 _1554_ (.A(_0110_),
    .B(_0112_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[27] ));
 sky130_fd_sc_hd__mux2i_2 _1555_ (.A0(net49),
    .A1(net111),
    .S(_0869_),
    .Y(_0113_));
 sky130_fd_sc_hd__nor3_1 _1556_ (.A(_0870_),
    .B(_0995_),
    .C(net24),
    .Y(_0114_));
 sky130_fd_sc_hd__a211oi_4 _1557_ (.A1(_0995_),
    .A2(_0113_),
    .B1(_0114_),
    .C1(_0884_),
    .Y(_0115_));
 sky130_fd_sc_hd__or3_1 _1558_ (.A(_0869_),
    .B(_0927_),
    .C(net80),
    .X(_0116_));
 sky130_fd_sc_hd__nand2b_1 _1559_ (.A_N(net24),
    .B(_0927_),
    .Y(_0117_));
 sky130_fd_sc_hd__a31o_1 _1560_ (.A1(_0884_),
    .A2(_0116_),
    .A3(_0117_),
    .B1(_0782_),
    .X(_0118_));
 sky130_fd_sc_hd__a21o_1 _1561_ (.A1(_0784_),
    .A2(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[28] ),
    .B1(_0771_),
    .X(_0119_));
 sky130_fd_sc_hd__nor2b_1 _1562_ (.A(net24),
    .B_N(_0884_),
    .Y(_0120_));
 sky130_fd_sc_hd__nor4_1 _1563_ (.A(_0883_),
    .B(_0995_),
    .C(_0853_),
    .D(net141),
    .Y(_0121_));
 sky130_fd_sc_hd__o211ai_2 _1564_ (.A1(_0120_),
    .A2(_0121_),
    .B1(_0771_),
    .C1(_0870_),
    .Y(_0122_));
 sky130_fd_sc_hd__o211ai_4 _1565_ (.A1(_0115_),
    .A2(_0118_),
    .B1(_0119_),
    .C1(_0122_),
    .Y(_0123_));
 sky130_fd_sc_hd__nand2_1 _1566_ (.A(_0110_),
    .B(_0111_),
    .Y(_0124_));
 sky130_fd_sc_hd__nor4_1 _1567_ (.A(_0970_),
    .B(_0076_),
    .C(_0077_),
    .D(_0124_),
    .Y(_0125_));
 sky130_fd_sc_hd__xnor2_1 _1568_ (.A(_0123_),
    .B(_0125_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[28] ));
 sky130_fd_sc_hd__mux2i_1 _1569_ (.A0(net50),
    .A1(net112),
    .S(_0870_),
    .Y(_0126_));
 sky130_fd_sc_hd__o2bb2ai_1 _1570_ (.A1_N(net142),
    .A2_N(_0031_),
    .B1(_0126_),
    .B2(_0868_),
    .Y(_0127_));
 sky130_fd_sc_hd__nand2_1 _1571_ (.A(_0884_),
    .B(net25),
    .Y(_0128_));
 sky130_fd_sc_hd__or4b_1 _1572_ (.A(_0900_),
    .B(_0869_),
    .C(_0927_),
    .D_N(net25),
    .X(_0129_));
 sky130_fd_sc_hd__o21ai_2 _1573_ (.A1(_0901_),
    .A2(_0128_),
    .B1(_0129_),
    .Y(_0130_));
 sky130_fd_sc_hd__nor4bb_1 _1574_ (.A(_0869_),
    .B(_0927_),
    .C_N(net81),
    .D_N(_0883_),
    .Y(_0131_));
 sky130_fd_sc_hd__nand2b_1 _1575_ (.A_N(_0131_),
    .B(_0914_),
    .Y(_0132_));
 sky130_fd_sc_hd__nor2b_1 _1576_ (.A(_0774_),
    .B_N(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[29] ),
    .Y(_0133_));
 sky130_fd_sc_hd__o32ai_4 _1577_ (.A1(_0127_),
    .A2(_0130_),
    .A3(_0132_),
    .B1(_0133_),
    .B2(_0899_),
    .Y(_0134_));
 sky130_fd_sc_hd__nor3_1 _1578_ (.A(_0102_),
    .B(_0109_),
    .C(_0123_),
    .Y(_0135_));
 sky130_fd_sc_hd__nand2_1 _1579_ (.A(_0111_),
    .B(_0135_),
    .Y(_0136_));
 sky130_fd_sc_hd__nor4_1 _1580_ (.A(_0984_),
    .B(_0076_),
    .C(_0077_),
    .D(_0136_),
    .Y(_0137_));
 sky130_fd_sc_hd__xnor2_1 _1581_ (.A(_0134_),
    .B(_0137_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[29] ));
 sky130_fd_sc_hd__mux2i_2 _1582_ (.A0(net26),
    .A1(net83),
    .S(_0901_),
    .Y(_0138_));
 sky130_fd_sc_hd__nand2_1 _1583_ (.A(_0924_),
    .B(net26),
    .Y(_0139_));
 sky130_fd_sc_hd__mux2_1 _1584_ (.A0(net52),
    .A1(net114),
    .S(_0870_),
    .X(_0140_));
 sky130_fd_sc_hd__a22oi_2 _1585_ (.A1(net143),
    .A2(_0031_),
    .B1(_0140_),
    .B2(_1051_),
    .Y(_0141_));
 sky130_fd_sc_hd__o221ai_4 _1586_ (.A1(_0924_),
    .A2(_0138_),
    .B1(_0139_),
    .B2(_0885_),
    .C1(_0141_),
    .Y(_0142_));
 sky130_fd_sc_hd__nand2_1 _1587_ (.A(_0784_),
    .B(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[30] ),
    .Y(_0143_));
 sky130_fd_sc_hd__nor2_1 _1588_ (.A(_0899_),
    .B(_0143_),
    .Y(_0144_));
 sky130_fd_sc_hd__a21oi_1 _1589_ (.A1(_0899_),
    .A2(_0142_),
    .B1(_0144_),
    .Y(_0145_));
 sky130_fd_sc_hd__nor4_1 _1590_ (.A(_0102_),
    .B(_0109_),
    .C(_0123_),
    .D(_0134_),
    .Y(_0146_));
 sky130_fd_sc_hd__nand2_1 _1591_ (.A(_0111_),
    .B(_0146_),
    .Y(_0147_));
 sky130_fd_sc_hd__nor4_1 _1592_ (.A(_0970_),
    .B(_0076_),
    .C(_0077_),
    .D(_0147_),
    .Y(_0148_));
 sky130_fd_sc_hd__xnor2_1 _1593_ (.A(_0145_),
    .B(_0148_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[30] ));
 sky130_fd_sc_hd__nor2b_1 _1594_ (.A(_0774_),
    .B_N(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[31] ),
    .Y(_0149_));
 sky130_fd_sc_hd__mux2i_1 _1595_ (.A0(net53),
    .A1(net115),
    .S(_0870_),
    .Y(_0150_));
 sky130_fd_sc_hd__nand2_1 _1596_ (.A(net144),
    .B(_0031_),
    .Y(_0151_));
 sky130_fd_sc_hd__o21ai_0 _1597_ (.A1(_0868_),
    .A2(_0150_),
    .B1(_0151_),
    .Y(_0152_));
 sky130_fd_sc_hd__a221oi_2 _1598_ (.A1(net84),
    .A2(_0855_),
    .B1(_1049_),
    .B2(net27),
    .C1(_0152_),
    .Y(_0153_));
 sky130_fd_sc_hd__nand2_1 _1599_ (.A(_0017_),
    .B(_0153_),
    .Y(_0154_));
 sky130_fd_sc_hd__o21ai_0 _1600_ (.A1(_0017_),
    .A2(_0149_),
    .B1(_0154_),
    .Y(_0155_));
 sky130_fd_sc_hd__nand3b_1 _1601_ (.A_N(_0145_),
    .B(_0146_),
    .C(_0111_),
    .Y(_0156_));
 sky130_fd_sc_hd__nor4_4 _1602_ (.A(_0984_),
    .B(_1023_),
    .C(_0057_),
    .D(_0156_),
    .Y(_0157_));
 sky130_fd_sc_hd__xnor2_1 _1603_ (.A(_0155_),
    .B(_0157_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[31] ));
 sky130_fd_sc_hd__nor2_1 _1604_ (.A(_0940_),
    .B(_0943_),
    .Y(_0158_));
 sky130_fd_sc_hd__nor2b_1 _1605_ (.A(_0158_),
    .B_N(_0945_),
    .Y(_0159_));
 sky130_fd_sc_hd__xor2_1 _1606_ (.A(_1068_),
    .B(_0159_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[4] ));
 sky130_fd_sc_hd__nand3_1 _1607_ (.A(_1066_),
    .B(_1067_),
    .C(_0159_),
    .Y(_0160_));
 sky130_fd_sc_hd__xor2_1 _1608_ (.A(_0958_),
    .B(_0160_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[5] ));
 sky130_fd_sc_hd__o21a_1 _1609_ (.A1(_0946_),
    .A2(_0958_),
    .B1(_0952_),
    .X(_0161_));
 sky130_fd_sc_hd__nor2_1 _1610_ (.A(_0959_),
    .B(_0161_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[6] ));
 sky130_fd_sc_hd__a21oi_1 _1611_ (.A1(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[7] ),
    .A2(_1033_),
    .B1(_0936_),
    .Y(_0162_));
 sky130_fd_sc_hd__xnor2_1 _1612_ (.A(_0982_),
    .B(_0162_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[7] ));
 sky130_fd_sc_hd__nor2b_1 _1613_ (.A(_0162_),
    .B_N(_0959_),
    .Y(_0163_));
 sky130_fd_sc_hd__nor2_2 _1614_ (.A(_0931_),
    .B(_0930_),
    .Y(_0164_));
 sky130_fd_sc_hd__a22oi_1 _1615_ (.A1(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[8] ),
    .A2(_1033_),
    .B1(_0164_),
    .B2(_0017_),
    .Y(_0165_));
 sky130_fd_sc_hd__xnor2_1 _1616_ (.A(_0163_),
    .B(_0165_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[8] ));
 sky130_fd_sc_hd__o21ai_0 _1617_ (.A1(_0937_),
    .A2(_0938_),
    .B1(_0982_),
    .Y(_0166_));
 sky130_fd_sc_hd__xnor2_1 _1618_ (.A(_0968_),
    .B(_0166_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[9] ));
 sky130_fd_sc_hd__nand2_8 _1619_ (.A(_1033_),
    .B(_0864_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ));
 sky130_fd_sc_hd__o2111ai_4 _1620_ (.A1(_0837_),
    .A2(_0840_),
    .B1(_0843_),
    .C1(_0768_),
    .D1(net154),
    .Y(_0167_));
 sky130_fd_sc_hd__or2_2 _1621_ (.A(_0841_),
    .B(_0167_),
    .X(_0168_));
 sky130_fd_sc_hd__nor2_2 _1622_ (.A(\gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0] ),
    .B(_0838_),
    .Y(_0169_));
 sky130_fd_sc_hd__xnor2_1 _1623_ (.A(_0839_),
    .B(_0167_),
    .Y(_0170_));
 sky130_fd_sc_hd__nand2_2 _1624_ (.A(_0169_),
    .B(_0170_),
    .Y(_0171_));
 sky130_fd_sc_hd__nand2_8 _1625_ (.A(_0168_),
    .B(_0171_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ));
 sky130_fd_sc_hd__inv_1 _1626_ (.A(_0167_),
    .Y(_0172_));
 sky130_fd_sc_hd__nand3_1 _1627_ (.A(_0877_),
    .B(_0841_),
    .C(_0167_),
    .Y(_0173_));
 sky130_fd_sc_hd__nand2_1 _1628_ (.A(_0168_),
    .B(_0173_),
    .Y(_0174_));
 sky130_fd_sc_hd__a22o_4 _1629_ (.A1(_0846_),
    .A2(_0172_),
    .B1(_0174_),
    .B2(_0169_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[1] ));
 sky130_fd_sc_hd__mux2_1 _1630_ (.A0(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1] ),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_d[2] ),
    .S(_0841_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_d[0] ));
 sky130_fd_sc_hd__mux2_1 _1631_ (.A0(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_d[2] ),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[2] ),
    .S(_0846_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_d[1] ));
 sky130_fd_sc_hd__buf_4 _1632_ (.A(_0017_),
    .X(_0175_));
 sky130_fd_sc_hd__nor2_1 _1633_ (.A(_0175_),
    .B(_1061_),
    .Y(_0176_));
 sky130_fd_sc_hd__mux2_1 _1634_ (.A0(net40),
    .A1(net102),
    .S(_0870_),
    .X(_0177_));
 sky130_fd_sc_hd__a221oi_4 _1635_ (.A1(net71),
    .A2(_0855_),
    .B1(_1051_),
    .B2(_0177_),
    .C1(_0880_),
    .Y(_0178_));
 sky130_fd_sc_hd__nor3_1 _1636_ (.A(_0834_),
    .B(_0176_),
    .C(_0178_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[1] ));
 sky130_fd_sc_hd__inv_1 _1637_ (.A(net348),
    .Y(_0179_));
 sky130_fd_sc_hd__and2_1 _1638_ (.A(_1058_),
    .B(net372),
    .X(_0180_));
 sky130_fd_sc_hd__and4_2 _1639_ (.A(net373),
    .B(net374),
    .C(net375),
    .D(net376),
    .X(_0181_));
 sky130_fd_sc_hd__nand4_4 _1640_ (.A(net377),
    .B(net378),
    .C(_0180_),
    .D(_0181_),
    .Y(_0182_));
 sky130_fd_sc_hd__o21ai_0 _1641_ (.A1(_0179_),
    .A2(_0182_),
    .B1(net349),
    .Y(_0183_));
 sky130_fd_sc_hd__or3_1 _1642_ (.A(_0179_),
    .B(net349),
    .C(_0182_),
    .X(_0184_));
 sky130_fd_sc_hd__a311oi_1 _1643_ (.A1(_0875_),
    .A2(_0183_),
    .A3(_0184_),
    .B1(_0834_),
    .C1(_0979_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[11] ));
 sky130_fd_sc_hd__nand3_2 _1644_ (.A(net377),
    .B(net378),
    .C(_0181_),
    .Y(_0185_));
 sky130_fd_sc_hd__a21o_1 _1645_ (.A1(_1056_),
    .A2(_1063_),
    .B1(_1062_),
    .X(_0186_));
 sky130_fd_sc_hd__nand2_2 _1646_ (.A(net372),
    .B(_0186_),
    .Y(_0187_));
 sky130_fd_sc_hd__nor2_1 _1647_ (.A(_0185_),
    .B(_0187_),
    .Y(_0188_));
 sky130_fd_sc_hd__nand3_1 _1648_ (.A(net348),
    .B(net349),
    .C(_0188_),
    .Y(_0189_));
 sky130_fd_sc_hd__xor2_1 _1649_ (.A(net350),
    .B(_0189_),
    .X(_0190_));
 sky130_fd_sc_hd__a21o_2 _1650_ (.A1(_0865_),
    .A2(_0994_),
    .B1(_0989_),
    .X(_0191_));
 sky130_fd_sc_hd__nor2_1 _1651_ (.A(_0875_),
    .B(_0191_),
    .Y(_0192_));
 sky130_fd_sc_hd__buf_4 _1652_ (.A(_0834_),
    .X(_0193_));
 sky130_fd_sc_hd__a211oi_1 _1653_ (.A1(_0881_),
    .A2(_0190_),
    .B1(_0192_),
    .C1(_0193_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[12] ));
 sky130_fd_sc_hd__nand3_1 _1654_ (.A(net348),
    .B(net349),
    .C(net350),
    .Y(_0194_));
 sky130_fd_sc_hd__nor2_1 _1655_ (.A(_0182_),
    .B(_0194_),
    .Y(_0195_));
 sky130_fd_sc_hd__xnor2_1 _1656_ (.A(net351),
    .B(_0195_),
    .Y(_0196_));
 sky130_fd_sc_hd__a21o_1 _1657_ (.A1(_0865_),
    .A2(_1008_),
    .B1(_1007_),
    .X(_0197_));
 sky130_fd_sc_hd__nor2_2 _1658_ (.A(_0880_),
    .B(_0197_),
    .Y(_0198_));
 sky130_fd_sc_hd__a211oi_1 _1659_ (.A1(_0881_),
    .A2(_0196_),
    .B1(_0198_),
    .C1(_0193_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[13] ));
 sky130_fd_sc_hd__nand4_4 _1660_ (.A(net348),
    .B(net349),
    .C(net350),
    .D(net351),
    .Y(_0199_));
 sky130_fd_sc_hd__nor3_1 _1661_ (.A(_0185_),
    .B(_0187_),
    .C(_0199_),
    .Y(_0200_));
 sky130_fd_sc_hd__xor2_1 _1662_ (.A(net352),
    .B(_0200_),
    .X(_0201_));
 sky130_fd_sc_hd__nor2_1 _1663_ (.A(_0044_),
    .B(_0201_),
    .Y(_0202_));
 sky130_fd_sc_hd__a211oi_1 _1664_ (.A1(_0175_),
    .A2(_1017_),
    .B1(_0202_),
    .C1(_0193_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[14] ));
 sky130_fd_sc_hd__nor2_1 _1665_ (.A(_0182_),
    .B(_0199_),
    .Y(_0203_));
 sky130_fd_sc_hd__nand2_1 _1666_ (.A(net352),
    .B(_0203_),
    .Y(_0204_));
 sky130_fd_sc_hd__xor2_1 _1667_ (.A(net353),
    .B(_0204_),
    .X(_0205_));
 sky130_fd_sc_hd__o21a_1 _1668_ (.A1(_0017_),
    .A2(_0205_),
    .B1(_1032_),
    .X(_0206_));
 sky130_fd_sc_hd__nor2_1 _1669_ (.A(_0835_),
    .B(_0206_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[15] ));
 sky130_fd_sc_hd__nand3_1 _1670_ (.A(net352),
    .B(net353),
    .C(_0200_),
    .Y(_0207_));
 sky130_fd_sc_hd__xnor2_1 _1671_ (.A(net354),
    .B(_0207_),
    .Y(_0208_));
 sky130_fd_sc_hd__a21oi_1 _1672_ (.A1(_0875_),
    .A2(_0208_),
    .B1(_1043_),
    .Y(_0209_));
 sky130_fd_sc_hd__nor2_1 _1673_ (.A(_0835_),
    .B(_0209_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[16] ));
 sky130_fd_sc_hd__nand4_1 _1674_ (.A(net352),
    .B(net353),
    .C(net354),
    .D(_0203_),
    .Y(_0210_));
 sky130_fd_sc_hd__xnor2_1 _1675_ (.A(net355),
    .B(_0210_),
    .Y(_0211_));
 sky130_fd_sc_hd__nor2_1 _1676_ (.A(_0044_),
    .B(_0211_),
    .Y(_0212_));
 sky130_fd_sc_hd__a211oi_1 _1677_ (.A1(_0175_),
    .A2(_1053_),
    .B1(_0212_),
    .C1(_0193_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[17] ));
 sky130_fd_sc_hd__nand4_4 _1678_ (.A(net352),
    .B(net353),
    .C(net354),
    .D(net355),
    .Y(_0213_));
 sky130_fd_sc_hd__nor4_4 _1679_ (.A(_0185_),
    .B(_0187_),
    .C(_0199_),
    .D(_0213_),
    .Y(_0214_));
 sky130_fd_sc_hd__xnor2_1 _1680_ (.A(net356),
    .B(_0214_),
    .Y(_0215_));
 sky130_fd_sc_hd__nor2_1 _1681_ (.A(_0880_),
    .B(_0009_),
    .Y(_0216_));
 sky130_fd_sc_hd__a211oi_1 _1682_ (.A1(_0881_),
    .A2(_0215_),
    .B1(_0216_),
    .C1(_0193_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[18] ));
 sky130_fd_sc_hd__nor3_1 _1683_ (.A(_0182_),
    .B(_0199_),
    .C(_0213_),
    .Y(_0217_));
 sky130_fd_sc_hd__nand2_1 _1684_ (.A(net356),
    .B(_0217_),
    .Y(_0218_));
 sky130_fd_sc_hd__xnor2_1 _1685_ (.A(net357),
    .B(_0218_),
    .Y(_0219_));
 sky130_fd_sc_hd__nor2_1 _1686_ (.A(_0044_),
    .B(_0219_),
    .Y(_0220_));
 sky130_fd_sc_hd__nor2_1 _1687_ (.A(_0875_),
    .B(_0016_),
    .Y(_0221_));
 sky130_fd_sc_hd__nor3_1 _1688_ (.A(_0834_),
    .B(_0220_),
    .C(_0221_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[19] ));
 sky130_fd_sc_hd__nand3_1 _1689_ (.A(net356),
    .B(net357),
    .C(_0214_),
    .Y(_0222_));
 sky130_fd_sc_hd__xor2_1 _1690_ (.A(net359),
    .B(_0222_),
    .X(_0223_));
 sky130_fd_sc_hd__nor2_1 _1691_ (.A(_0880_),
    .B(_0026_),
    .Y(_0224_));
 sky130_fd_sc_hd__a211oi_1 _1692_ (.A1(_0881_),
    .A2(_0223_),
    .B1(_0224_),
    .C1(_0193_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[20] ));
 sky130_fd_sc_hd__nor2_1 _1693_ (.A(_0044_),
    .B(_1059_),
    .Y(_0225_));
 sky130_fd_sc_hd__a211oi_1 _1694_ (.A1(_0175_),
    .A2(_0873_),
    .B1(_0225_),
    .C1(_0193_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[2] ));
 sky130_fd_sc_hd__and3_1 _1695_ (.A(net356),
    .B(net357),
    .C(net359),
    .X(_0226_));
 sky130_fd_sc_hd__nand2_1 _1696_ (.A(_0217_),
    .B(_0226_),
    .Y(_0227_));
 sky130_fd_sc_hd__xor2_1 _1697_ (.A(net360),
    .B(_0227_),
    .X(_0228_));
 sky130_fd_sc_hd__o21a_1 _1698_ (.A1(_0017_),
    .A2(_0228_),
    .B1(_0038_),
    .X(_0229_));
 sky130_fd_sc_hd__nor2_1 _1699_ (.A(_0835_),
    .B(_0229_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[21] ));
 sky130_fd_sc_hd__nand3_1 _1700_ (.A(net360),
    .B(_0214_),
    .C(_0226_),
    .Y(_0230_));
 sky130_fd_sc_hd__xor2_1 _1701_ (.A(net361),
    .B(_0230_),
    .X(_0231_));
 sky130_fd_sc_hd__a211oi_1 _1702_ (.A1(_0881_),
    .A2(_0231_),
    .B1(_0051_),
    .C1(_0193_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[22] ));
 sky130_fd_sc_hd__and3_1 _1703_ (.A(net360),
    .B(net361),
    .C(_0226_),
    .X(_0232_));
 sky130_fd_sc_hd__nor4b_4 _1704_ (.A(_0182_),
    .B(_0199_),
    .C(_0213_),
    .D_N(_0232_),
    .Y(_0233_));
 sky130_fd_sc_hd__xor2_1 _1705_ (.A(net362),
    .B(_0233_),
    .X(_0234_));
 sky130_fd_sc_hd__a21boi_0 _1706_ (.A1(_0875_),
    .A2(_0234_),
    .B1_N(_0064_),
    .Y(_0235_));
 sky130_fd_sc_hd__nor2_1 _1707_ (.A(_0835_),
    .B(_0235_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[23] ));
 sky130_fd_sc_hd__o21ai_4 _1708_ (.A1(_0995_),
    .A2(_0072_),
    .B1(_0071_),
    .Y(_0236_));
 sky130_fd_sc_hd__nand3_1 _1709_ (.A(net362),
    .B(_0214_),
    .C(_0232_),
    .Y(_0237_));
 sky130_fd_sc_hd__xnor2_1 _1710_ (.A(net363),
    .B(_0237_),
    .Y(_0238_));
 sky130_fd_sc_hd__mux2i_1 _1711_ (.A0(_0236_),
    .A1(_0238_),
    .S(_0875_),
    .Y(_0239_));
 sky130_fd_sc_hd__nor2_1 _1712_ (.A(_0835_),
    .B(_0239_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[24] ));
 sky130_fd_sc_hd__nand3_1 _1713_ (.A(_0884_),
    .B(_0082_),
    .C(_0083_),
    .Y(_0240_));
 sky130_fd_sc_hd__a21oi_1 _1714_ (.A1(_0086_),
    .A2(_0087_),
    .B1(_0926_),
    .Y(_0241_));
 sky130_fd_sc_hd__a21o_2 _1715_ (.A1(_0081_),
    .A2(_0240_),
    .B1(_0241_),
    .X(_0242_));
 sky130_fd_sc_hd__nand3_1 _1716_ (.A(net362),
    .B(net363),
    .C(_0233_),
    .Y(_0243_));
 sky130_fd_sc_hd__xnor2_1 _1717_ (.A(net364),
    .B(_0243_),
    .Y(_0244_));
 sky130_fd_sc_hd__nor2_1 _1718_ (.A(_0044_),
    .B(_0244_),
    .Y(_0245_));
 sky130_fd_sc_hd__a211oi_1 _1719_ (.A1(_0175_),
    .A2(_0242_),
    .B1(_0245_),
    .C1(_0193_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[25] ));
 sky130_fd_sc_hd__and3_1 _1720_ (.A(net362),
    .B(net363),
    .C(net364),
    .X(_0246_));
 sky130_fd_sc_hd__nand3_1 _1721_ (.A(_0214_),
    .B(_0232_),
    .C(_0246_),
    .Y(_0247_));
 sky130_fd_sc_hd__xor2_1 _1722_ (.A(net365),
    .B(_0247_),
    .X(_0248_));
 sky130_fd_sc_hd__a21o_1 _1723_ (.A1(_0865_),
    .A2(_0096_),
    .B1(_0095_),
    .X(_0249_));
 sky130_fd_sc_hd__nor2_2 _1724_ (.A(_0880_),
    .B(_0249_),
    .Y(_0250_));
 sky130_fd_sc_hd__a211oi_1 _1725_ (.A1(_0881_),
    .A2(_0248_),
    .B1(_0250_),
    .C1(_0193_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[26] ));
 sky130_fd_sc_hd__and2_0 _1726_ (.A(net365),
    .B(_0246_),
    .X(_0251_));
 sky130_fd_sc_hd__nand2_1 _1727_ (.A(_0233_),
    .B(_0251_),
    .Y(_0252_));
 sky130_fd_sc_hd__xor2_1 _1728_ (.A(net366),
    .B(_0252_),
    .X(_0253_));
 sky130_fd_sc_hd__a211oi_1 _1729_ (.A1(_0881_),
    .A2(_0253_),
    .B1(_0109_),
    .C1(_0834_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[27] ));
 sky130_fd_sc_hd__and3_1 _1730_ (.A(_0884_),
    .B(_0116_),
    .C(_0117_),
    .X(_0254_));
 sky130_fd_sc_hd__o21ai_1 _1731_ (.A1(_0120_),
    .A2(_0121_),
    .B1(_0870_),
    .Y(_0255_));
 sky130_fd_sc_hd__o21ai_4 _1732_ (.A1(_0115_),
    .A2(_0254_),
    .B1(_0255_),
    .Y(_0256_));
 sky130_fd_sc_hd__nand4_1 _1733_ (.A(net366),
    .B(_0214_),
    .C(_0232_),
    .D(_0251_),
    .Y(_0257_));
 sky130_fd_sc_hd__xnor2_1 _1734_ (.A(net367),
    .B(_0257_),
    .Y(_0258_));
 sky130_fd_sc_hd__nor2_1 _1735_ (.A(_0044_),
    .B(_0258_),
    .Y(_0259_));
 sky130_fd_sc_hd__a211oi_1 _1736_ (.A1(_0175_),
    .A2(_0256_),
    .B1(_0259_),
    .C1(_0834_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[28] ));
 sky130_fd_sc_hd__or3_4 _1737_ (.A(_0127_),
    .B(_0130_),
    .C(_0131_),
    .X(_0260_));
 sky130_fd_sc_hd__and3_1 _1738_ (.A(net366),
    .B(net367),
    .C(_0251_),
    .X(_0261_));
 sky130_fd_sc_hd__nand2_1 _1739_ (.A(_0233_),
    .B(_0261_),
    .Y(_0262_));
 sky130_fd_sc_hd__xnor2_1 _1740_ (.A(net368),
    .B(_0262_),
    .Y(_0263_));
 sky130_fd_sc_hd__mux2i_1 _1741_ (.A0(_0260_),
    .A1(_0263_),
    .S(_0875_),
    .Y(_0264_));
 sky130_fd_sc_hd__nor2_1 _1742_ (.A(_0835_),
    .B(_0264_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[29] ));
 sky130_fd_sc_hd__nand4_1 _1743_ (.A(net368),
    .B(_0214_),
    .C(_0232_),
    .D(_0261_),
    .Y(_0265_));
 sky130_fd_sc_hd__xor2_1 _1744_ (.A(net370),
    .B(_0265_),
    .X(_0266_));
 sky130_fd_sc_hd__buf_6 _1745_ (.A(_0784_),
    .X(_0267_));
 sky130_fd_sc_hd__nand3_1 _1746_ (.A(_0175_),
    .B(_0267_),
    .C(_0142_),
    .Y(_0268_));
 sky130_fd_sc_hd__o21ai_0 _1747_ (.A1(_0785_),
    .A2(_0266_),
    .B1(_0268_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[30] ));
 sky130_fd_sc_hd__xnor2_1 _1748_ (.A(_1058_),
    .B(net372),
    .Y(_0269_));
 sky130_fd_sc_hd__a221oi_1 _1749_ (.A1(_0856_),
    .A2(_0861_),
    .B1(_0269_),
    .B2(_0875_),
    .C1(_0834_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[3] ));
 sky130_fd_sc_hd__nand4_1 _1750_ (.A(net368),
    .B(net370),
    .C(_0233_),
    .D(_0261_),
    .Y(_0270_));
 sky130_fd_sc_hd__xnor2_1 _1751_ (.A(net371),
    .B(_0270_),
    .Y(_0271_));
 sky130_fd_sc_hd__o211a_1 _1752_ (.A1(_0175_),
    .A2(_0271_),
    .B1(_0154_),
    .C1(_0267_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[31] ));
 sky130_fd_sc_hd__xor2_1 _1753_ (.A(net373),
    .B(_0187_),
    .X(_0272_));
 sky130_fd_sc_hd__a211oi_1 _1754_ (.A1(_0881_),
    .A2(_0272_),
    .B1(_0158_),
    .C1(_0834_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[4] ));
 sky130_fd_sc_hd__nand2_1 _1755_ (.A(net373),
    .B(_0180_),
    .Y(_0273_));
 sky130_fd_sc_hd__xnor2_1 _1756_ (.A(net374),
    .B(_0273_),
    .Y(_0274_));
 sky130_fd_sc_hd__o22ai_1 _1757_ (.A1(_0957_),
    .A2(_0955_),
    .B1(_0274_),
    .B2(_0175_),
    .Y(_0275_));
 sky130_fd_sc_hd__nor2_1 _1758_ (.A(_0835_),
    .B(_0275_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[5] ));
 sky130_fd_sc_hd__nand2_1 _1759_ (.A(net373),
    .B(net374),
    .Y(_0276_));
 sky130_fd_sc_hd__nor2_1 _1760_ (.A(_0276_),
    .B(_0187_),
    .Y(_0277_));
 sky130_fd_sc_hd__xor2_1 _1761_ (.A(net375),
    .B(_0277_),
    .X(_0278_));
 sky130_fd_sc_hd__o221a_1 _1762_ (.A1(_0951_),
    .A2(_0949_),
    .B1(_0278_),
    .B2(_0044_),
    .C1(_0267_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[6] ));
 sky130_fd_sc_hd__nand4_1 _1763_ (.A(net373),
    .B(net374),
    .C(net375),
    .D(_0180_),
    .Y(_0279_));
 sky130_fd_sc_hd__xor2_1 _1764_ (.A(net376),
    .B(_0279_),
    .X(_0280_));
 sky130_fd_sc_hd__nor2_1 _1765_ (.A(_0044_),
    .B(_0280_),
    .Y(_0281_));
 sky130_fd_sc_hd__nor2_1 _1766_ (.A(_0936_),
    .B(_0281_),
    .Y(_0282_));
 sky130_fd_sc_hd__nor2_1 _1767_ (.A(_0835_),
    .B(_0282_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[7] ));
 sky130_fd_sc_hd__nand3_1 _1768_ (.A(net372),
    .B(_0181_),
    .C(_0186_),
    .Y(_0283_));
 sky130_fd_sc_hd__xnor2_1 _1769_ (.A(net377),
    .B(_0283_),
    .Y(_0284_));
 sky130_fd_sc_hd__o21ai_1 _1770_ (.A1(_0931_),
    .A2(_0930_),
    .B1(_0044_),
    .Y(_0285_));
 sky130_fd_sc_hd__o211a_1 _1771_ (.A1(_0175_),
    .A2(_0284_),
    .B1(_0285_),
    .C1(_0267_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[8] ));
 sky130_fd_sc_hd__nand3_1 _1772_ (.A(net377),
    .B(_0180_),
    .C(_0181_),
    .Y(_0286_));
 sky130_fd_sc_hd__xnor2_1 _1773_ (.A(net378),
    .B(_0286_),
    .Y(_0287_));
 sky130_fd_sc_hd__nor2_1 _1774_ (.A(_0965_),
    .B(_0966_),
    .Y(_0288_));
 sky130_fd_sc_hd__a21oi_1 _1775_ (.A1(_0875_),
    .A2(_0287_),
    .B1(_0288_),
    .Y(_0289_));
 sky130_fd_sc_hd__nor2_1 _1776_ (.A(_0835_),
    .B(_0289_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[9] ));
 sky130_fd_sc_hd__xnor2_1 _1777_ (.A(net348),
    .B(_0188_),
    .Y(_0290_));
 sky130_fd_sc_hd__nor2_2 _1778_ (.A(_0880_),
    .B(_0913_),
    .Y(_0291_));
 sky130_fd_sc_hd__a211oi_1 _1779_ (.A1(_0881_),
    .A2(_0290_),
    .B1(_0291_),
    .C1(_0834_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[10] ));
 sky130_fd_sc_hd__nand2_8 _1780_ (.A(_1033_),
    .B(_0844_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_en ));
 sky130_fd_sc_hd__mux2i_2 _1781_ (.A0(net158),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[32] ),
    .S(\gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .Y(_0292_));
 sky130_fd_sc_hd__inv_1 _1782_ (.A(_0292_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[0] ));
 sky130_fd_sc_hd__mux2_1 _1783_ (.A0(net165),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[48] ),
    .S(_0876_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[16] ));
 sky130_fd_sc_hd__mux2_1 _1784_ (.A0(net166),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[49] ),
    .S(_0876_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[17] ));
 sky130_fd_sc_hd__mux2_1 _1785_ (.A0(net167),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[50] ),
    .S(_0876_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[18] ));
 sky130_fd_sc_hd__mux2_1 _1786_ (.A0(net168),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[51] ),
    .S(_0876_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[19] ));
 sky130_fd_sc_hd__mux2_1 _1787_ (.A0(net169),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[33] ),
    .S(_0776_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[1] ));
 sky130_fd_sc_hd__mux2_1 _1788_ (.A0(net170),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[52] ),
    .S(_0876_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[20] ));
 sky130_fd_sc_hd__mux2_1 _1789_ (.A0(net171),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[53] ),
    .S(_0876_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[21] ));
 sky130_fd_sc_hd__clkbuf_8 _1790_ (.A(_0821_),
    .X(_0293_));
 sky130_fd_sc_hd__mux2_1 _1791_ (.A0(net172),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[54] ),
    .S(_0293_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[22] ));
 sky130_fd_sc_hd__mux2_1 _1792_ (.A0(net173),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[55] ),
    .S(_0293_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[23] ));
 sky130_fd_sc_hd__mux2_1 _1793_ (.A0(net174),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[56] ),
    .S(_0293_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[24] ));
 sky130_fd_sc_hd__mux2_1 _1794_ (.A0(net175),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[57] ),
    .S(_0293_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[25] ));
 sky130_fd_sc_hd__mux2_1 _1795_ (.A0(net176),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[58] ),
    .S(_0293_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[26] ));
 sky130_fd_sc_hd__mux2_1 _1796_ (.A0(net177),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[59] ),
    .S(_0293_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[27] ));
 sky130_fd_sc_hd__mux2_1 _1797_ (.A0(net178),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[60] ),
    .S(_0293_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[28] ));
 sky130_fd_sc_hd__mux2_1 _1798_ (.A0(net179),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[61] ),
    .S(_0293_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[29] ));
 sky130_fd_sc_hd__mux2i_1 _1799_ (.A0(net180),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[34] ),
    .S(_0776_),
    .Y(_0294_));
 sky130_fd_sc_hd__inv_1 _1800_ (.A(_0294_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[2] ));
 sky130_fd_sc_hd__mux2_1 _1801_ (.A0(net181),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[62] ),
    .S(_0293_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[30] ));
 sky130_fd_sc_hd__mux2_1 _1802_ (.A0(net182),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[63] ),
    .S(_0293_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[31] ));
 sky130_fd_sc_hd__mux2_1 _1803_ (.A0(net158),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[64] ),
    .S(_0846_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[32] ));
 sky130_fd_sc_hd__mux2_1 _1804_ (.A0(net169),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[65] ),
    .S(_0846_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[33] ));
 sky130_fd_sc_hd__mux2_1 _1805_ (.A0(net180),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[66] ),
    .S(_0846_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[34] ));
 sky130_fd_sc_hd__mux2_1 _1806_ (.A0(net183),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[67] ),
    .S(_0846_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[35] ));
 sky130_fd_sc_hd__mux2_1 _1807_ (.A0(net184),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[68] ),
    .S(_0846_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[36] ));
 sky130_fd_sc_hd__clkbuf_8 _1808_ (.A(_0845_),
    .X(_0295_));
 sky130_fd_sc_hd__mux2_1 _1809_ (.A0(net185),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[69] ),
    .S(_0295_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[37] ));
 sky130_fd_sc_hd__mux2_1 _1810_ (.A0(net186),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[70] ),
    .S(_0295_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[38] ));
 sky130_fd_sc_hd__mux2_1 _1811_ (.A0(net187),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[71] ),
    .S(_0295_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[39] ));
 sky130_fd_sc_hd__mux2_1 _1812_ (.A0(net188),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[72] ),
    .S(_0295_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[40] ));
 sky130_fd_sc_hd__mux2_1 _1813_ (.A0(net189),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[73] ),
    .S(_0295_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[41] ));
 sky130_fd_sc_hd__mux2_1 _1814_ (.A0(net159),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[74] ),
    .S(_0295_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[42] ));
 sky130_fd_sc_hd__mux2_1 _1815_ (.A0(net160),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[75] ),
    .S(_0295_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[43] ));
 sky130_fd_sc_hd__mux2_1 _1816_ (.A0(net161),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[76] ),
    .S(_0295_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[44] ));
 sky130_fd_sc_hd__mux2_1 _1817_ (.A0(net162),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[77] ),
    .S(_0295_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[45] ));
 sky130_fd_sc_hd__mux2_1 _1818_ (.A0(net163),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[78] ),
    .S(_0295_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[46] ));
 sky130_fd_sc_hd__clkbuf_8 _1819_ (.A(_0845_),
    .X(_0296_));
 sky130_fd_sc_hd__mux2_1 _1820_ (.A0(net164),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[79] ),
    .S(_0296_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[47] ));
 sky130_fd_sc_hd__mux2_1 _1821_ (.A0(net165),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[80] ),
    .S(_0296_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[48] ));
 sky130_fd_sc_hd__mux2_1 _1822_ (.A0(net166),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[81] ),
    .S(_0296_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[49] ));
 sky130_fd_sc_hd__mux2_1 _1823_ (.A0(net167),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[82] ),
    .S(_0296_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[50] ));
 sky130_fd_sc_hd__mux2_1 _1824_ (.A0(net168),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[83] ),
    .S(_0296_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[51] ));
 sky130_fd_sc_hd__mux2_1 _1825_ (.A0(net170),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[84] ),
    .S(_0296_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[52] ));
 sky130_fd_sc_hd__mux2_1 _1826_ (.A0(net171),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[85] ),
    .S(_0296_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[53] ));
 sky130_fd_sc_hd__mux2_1 _1827_ (.A0(net172),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[86] ),
    .S(_0296_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[54] ));
 sky130_fd_sc_hd__mux2_1 _1828_ (.A0(net173),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[87] ),
    .S(_0296_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[55] ));
 sky130_fd_sc_hd__mux2_1 _1829_ (.A0(net174),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[88] ),
    .S(_0296_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[56] ));
 sky130_fd_sc_hd__mux2_1 _1830_ (.A0(net175),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[89] ),
    .S(_0845_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[57] ));
 sky130_fd_sc_hd__mux2_1 _1831_ (.A0(net176),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[90] ),
    .S(_0845_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[58] ));
 sky130_fd_sc_hd__mux2_1 _1832_ (.A0(net177),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[91] ),
    .S(_0845_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[59] ));
 sky130_fd_sc_hd__mux2_1 _1833_ (.A0(net178),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[92] ),
    .S(_0845_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[60] ));
 sky130_fd_sc_hd__mux2_1 _1834_ (.A0(net179),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[93] ),
    .S(_0845_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[61] ));
 sky130_fd_sc_hd__mux2_1 _1835_ (.A0(net181),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[94] ),
    .S(_0845_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[62] ));
 sky130_fd_sc_hd__mux2_1 _1836_ (.A0(net182),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[95] ),
    .S(_0845_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[63] ));
 sky130_fd_sc_hd__nand2_1 _1837_ (.A(_0169_),
    .B(_0167_),
    .Y(_0297_));
 sky130_fd_sc_hd__nor3_1 _1838_ (.A(_0821_),
    .B(_0169_),
    .C(_0167_),
    .Y(_0298_));
 sky130_fd_sc_hd__a311oi_1 _1839_ (.A1(_0839_),
    .A2(_0168_),
    .A3(_0297_),
    .B1(_0298_),
    .C1(_0785_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[0] ));
 sky130_fd_sc_hd__nand2_1 _1840_ (.A(_0846_),
    .B(_0172_),
    .Y(_0299_));
 sky130_fd_sc_hd__o21ai_0 _1841_ (.A1(_0169_),
    .A2(_0167_),
    .B1(_0876_),
    .Y(_0300_));
 sky130_fd_sc_hd__nand3_1 _1842_ (.A(_0877_),
    .B(_0169_),
    .C(_0167_),
    .Y(_0301_));
 sky130_fd_sc_hd__a31oi_1 _1843_ (.A1(_0299_),
    .A2(_0300_),
    .A3(_0301_),
    .B1(_0785_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[1] ));
 sky130_fd_sc_hd__a21oi_1 _1844_ (.A1(_0876_),
    .A2(_0169_),
    .B1(_0846_),
    .Y(_0302_));
 sky130_fd_sc_hd__nor3_1 _1845_ (.A(_0785_),
    .B(_0172_),
    .C(_0302_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[2] ));
 sky130_fd_sc_hd__buf_4 _1846_ (.A(_0769_),
    .X(_0303_));
 sky130_fd_sc_hd__buf_6 _1847_ (.A(_0772_),
    .X(_0304_));
 sky130_fd_sc_hd__buf_4 _1848_ (.A(_0772_),
    .X(_0305_));
 sky130_fd_sc_hd__nor2_1 _1849_ (.A(_0305_),
    .B(_0915_),
    .Y(_0306_));
 sky130_fd_sc_hd__a21oi_2 _1850_ (.A1(_0304_),
    .A2(_0913_),
    .B1(_0306_),
    .Y(_0307_));
 sky130_fd_sc_hd__buf_8 _1851_ (.A(_0769_),
    .X(_0308_));
 sky130_fd_sc_hd__clkbuf_4 _1852_ (.A(_0308_),
    .X(_0309_));
 sky130_fd_sc_hd__nand2_1 _1853_ (.A(_0309_),
    .B(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[10] ),
    .Y(_0310_));
 sky130_fd_sc_hd__o21ai_2 _1854_ (.A1(_0303_),
    .A2(_0307_),
    .B1(_0310_),
    .Y(net201));
 sky130_fd_sc_hd__a21oi_2 _1855_ (.A1(_0926_),
    .A2(_0975_),
    .B1(_0978_),
    .Y(_0311_));
 sky130_fd_sc_hd__mux2_1 _1856_ (.A0(_0311_),
    .A1(_0971_),
    .S(_0773_),
    .X(_0312_));
 sky130_fd_sc_hd__nand2_1 _1857_ (.A(_0309_),
    .B(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[11] ),
    .Y(_0313_));
 sky130_fd_sc_hd__o21ai_2 _1858_ (.A1(_0303_),
    .A2(_0312_),
    .B1(_0313_),
    .Y(net202));
 sky130_fd_sc_hd__buf_6 _1859_ (.A(_0769_),
    .X(_0314_));
 sky130_fd_sc_hd__nor2_1 _1860_ (.A(_0305_),
    .B(_0997_),
    .Y(_0315_));
 sky130_fd_sc_hd__a21oi_2 _1861_ (.A1(_0304_),
    .A2(_0191_),
    .B1(_0315_),
    .Y(_0316_));
 sky130_fd_sc_hd__nand2_1 _1862_ (.A(_0309_),
    .B(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[12] ),
    .Y(_0317_));
 sky130_fd_sc_hd__o21ai_2 _1863_ (.A1(_0314_),
    .A2(_0316_),
    .B1(_0317_),
    .Y(net203));
 sky130_fd_sc_hd__nor2_1 _1864_ (.A(_0305_),
    .B(_1009_),
    .Y(_0318_));
 sky130_fd_sc_hd__a21oi_2 _1865_ (.A1(_0304_),
    .A2(_0197_),
    .B1(_0318_),
    .Y(_0319_));
 sky130_fd_sc_hd__nand2_1 _1866_ (.A(_0309_),
    .B(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[13] ),
    .Y(_0320_));
 sky130_fd_sc_hd__o21ai_2 _1867_ (.A1(_0314_),
    .A2(_0319_),
    .B1(_0320_),
    .Y(net204));
 sky130_fd_sc_hd__buf_6 _1868_ (.A(_0773_),
    .X(_0321_));
 sky130_fd_sc_hd__clkbuf_8 _1869_ (.A(_0773_),
    .X(_0322_));
 sky130_fd_sc_hd__nor2_1 _1870_ (.A(_0322_),
    .B(_1017_),
    .Y(_0323_));
 sky130_fd_sc_hd__a31oi_2 _1871_ (.A1(_0267_),
    .A2(_0321_),
    .A3(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[14] ),
    .B1(_0323_),
    .Y(_0324_));
 sky130_fd_sc_hd__nand2_1 _1872_ (.A(_0309_),
    .B(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[14] ),
    .Y(_0325_));
 sky130_fd_sc_hd__o21ai_2 _1873_ (.A1(_0314_),
    .A2(_0324_),
    .B1(_0325_),
    .Y(net205));
 sky130_fd_sc_hd__or4_2 _1874_ (.A(_1027_),
    .B(_1028_),
    .C(_1029_),
    .D(_1031_),
    .X(_0326_));
 sky130_fd_sc_hd__nor2_4 _1875_ (.A(_0774_),
    .B(_0772_),
    .Y(_0327_));
 sky130_fd_sc_hd__a22oi_2 _1876_ (.A1(_0305_),
    .A2(_0326_),
    .B1(_0327_),
    .B2(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[15] ),
    .Y(_0328_));
 sky130_fd_sc_hd__nand2_1 _1877_ (.A(_0309_),
    .B(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[15] ),
    .Y(_0329_));
 sky130_fd_sc_hd__o21ai_2 _1878_ (.A1(_0314_),
    .A2(_0328_),
    .B1(_0329_),
    .Y(net206));
 sky130_fd_sc_hd__a2bb2oi_1 _1879_ (.A1_N(_0321_),
    .A2_N(_1042_),
    .B1(_0327_),
    .B2(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[16] ),
    .Y(_0330_));
 sky130_fd_sc_hd__nand2_1 _1880_ (.A(_0309_),
    .B(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[16] ),
    .Y(_0331_));
 sky130_fd_sc_hd__o21ai_2 _1881_ (.A1(_0314_),
    .A2(_0330_),
    .B1(_0331_),
    .Y(net207));
 sky130_fd_sc_hd__mux2_1 _1882_ (.A0(net8),
    .A1(_1054_),
    .S(_0773_),
    .X(_0332_));
 sky130_fd_sc_hd__nand2_1 _1883_ (.A(_0309_),
    .B(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[17] ),
    .Y(_0333_));
 sky130_fd_sc_hd__o21ai_2 _1884_ (.A1(_0314_),
    .A2(_0332_),
    .B1(_0333_),
    .Y(net208));
 sky130_fd_sc_hd__nor2_1 _1885_ (.A(_0772_),
    .B(_0010_),
    .Y(_0334_));
 sky130_fd_sc_hd__a21oi_1 _1886_ (.A1(_0304_),
    .A2(_0009_),
    .B1(_0334_),
    .Y(_0335_));
 sky130_fd_sc_hd__clkbuf_4 _1887_ (.A(_0308_),
    .X(_0336_));
 sky130_fd_sc_hd__nand2_1 _1888_ (.A(_0336_),
    .B(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[18] ),
    .Y(_0337_));
 sky130_fd_sc_hd__o21ai_2 _1889_ (.A1(_0314_),
    .A2(_0335_),
    .B1(_0337_),
    .Y(net209));
 sky130_fd_sc_hd__a22oi_1 _1890_ (.A1(_0305_),
    .A2(_0016_),
    .B1(_0327_),
    .B2(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[19] ),
    .Y(_0338_));
 sky130_fd_sc_hd__nand2_1 _1891_ (.A(_0336_),
    .B(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[19] ),
    .Y(_0339_));
 sky130_fd_sc_hd__o21ai_1 _1892_ (.A1(_0314_),
    .A2(_0338_),
    .B1(_0339_),
    .Y(net210));
 sky130_fd_sc_hd__a22oi_1 _1893_ (.A1(_0305_),
    .A2(_0026_),
    .B1(_0327_),
    .B2(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[20] ),
    .Y(_0340_));
 sky130_fd_sc_hd__nand2_1 _1894_ (.A(_0336_),
    .B(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[20] ),
    .Y(_0341_));
 sky130_fd_sc_hd__o21ai_1 _1895_ (.A1(_0314_),
    .A2(_0340_),
    .B1(_0341_),
    .Y(net211));
 sky130_fd_sc_hd__o21ai_2 _1896_ (.A1(_0033_),
    .A2(_0037_),
    .B1(_0772_),
    .Y(_0342_));
 sky130_fd_sc_hd__nand2_1 _1897_ (.A(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[21] ),
    .B(_0327_),
    .Y(_0343_));
 sky130_fd_sc_hd__a21oi_1 _1898_ (.A1(_0342_),
    .A2(_0343_),
    .B1(_0308_),
    .Y(_0344_));
 sky130_fd_sc_hd__a21o_1 _1899_ (.A1(_0303_),
    .A2(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[21] ),
    .B1(_0344_),
    .X(net212));
 sky130_fd_sc_hd__nor2_1 _1900_ (.A(_0321_),
    .B(_0050_),
    .Y(_0345_));
 sky130_fd_sc_hd__a21oi_1 _1901_ (.A1(_0321_),
    .A2(_0045_),
    .B1(_0345_),
    .Y(_0346_));
 sky130_fd_sc_hd__nand2_1 _1902_ (.A(_0336_),
    .B(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[22] ),
    .Y(_0347_));
 sky130_fd_sc_hd__o21ai_1 _1903_ (.A1(_0314_),
    .A2(_0346_),
    .B1(_0347_),
    .Y(net213));
 sky130_fd_sc_hd__o311ai_1 _1904_ (.A1(_0910_),
    .A2(_0060_),
    .A3(_0062_),
    .B1(_0063_),
    .C1(_0772_),
    .Y(_0348_));
 sky130_fd_sc_hd__nand3_1 _1905_ (.A(_0267_),
    .B(_0322_),
    .C(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[23] ),
    .Y(_0349_));
 sky130_fd_sc_hd__a21oi_1 _1906_ (.A1(_0348_),
    .A2(_0349_),
    .B1(_0308_),
    .Y(_0350_));
 sky130_fd_sc_hd__a21o_2 _1907_ (.A1(_0303_),
    .A2(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[23] ),
    .B1(_0350_),
    .X(net214));
 sky130_fd_sc_hd__buf_8 _1908_ (.A(_0769_),
    .X(_0351_));
 sky130_fd_sc_hd__and3_1 _1909_ (.A(_0267_),
    .B(_0322_),
    .C(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[24] ),
    .X(_0352_));
 sky130_fd_sc_hd__a21oi_2 _1910_ (.A1(_0304_),
    .A2(_0236_),
    .B1(_0352_),
    .Y(_0353_));
 sky130_fd_sc_hd__nand2_1 _1911_ (.A(_0336_),
    .B(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[24] ),
    .Y(_0354_));
 sky130_fd_sc_hd__o21ai_2 _1912_ (.A1(_0351_),
    .A2(_0353_),
    .B1(_0354_),
    .Y(net215));
 sky130_fd_sc_hd__nor2_1 _1913_ (.A(_0322_),
    .B(_0242_),
    .Y(_0355_));
 sky130_fd_sc_hd__a31oi_4 _1914_ (.A1(_0267_),
    .A2(_0321_),
    .A3(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[25] ),
    .B1(_0355_),
    .Y(_0356_));
 sky130_fd_sc_hd__nand2_1 _1915_ (.A(_0336_),
    .B(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[25] ),
    .Y(_0357_));
 sky130_fd_sc_hd__o21ai_2 _1916_ (.A1(_0351_),
    .A2(_0356_),
    .B1(_0357_),
    .Y(net216));
 sky130_fd_sc_hd__nor2_1 _1917_ (.A(_0772_),
    .B(_0097_),
    .Y(_0358_));
 sky130_fd_sc_hd__a21oi_2 _1918_ (.A1(_0304_),
    .A2(_0249_),
    .B1(_0358_),
    .Y(_0359_));
 sky130_fd_sc_hd__nand2_1 _1919_ (.A(_0336_),
    .B(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[26] ),
    .Y(_0360_));
 sky130_fd_sc_hd__o21ai_2 _1920_ (.A1(_0351_),
    .A2(_0359_),
    .B1(_0360_),
    .Y(net217));
 sky130_fd_sc_hd__inv_1 _1921_ (.A(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[27] ),
    .Y(_0361_));
 sky130_fd_sc_hd__a21oi_1 _1922_ (.A1(_0926_),
    .A2(_0105_),
    .B1(_0108_),
    .Y(_0362_));
 sky130_fd_sc_hd__nor2_1 _1923_ (.A(_0321_),
    .B(_0362_),
    .Y(_0363_));
 sky130_fd_sc_hd__a311oi_4 _1924_ (.A1(_0267_),
    .A2(_0321_),
    .A3(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[27] ),
    .B1(_0308_),
    .C1(_0363_),
    .Y(_0364_));
 sky130_fd_sc_hd__a21oi_2 _1925_ (.A1(_0309_),
    .A2(_0361_),
    .B1(_0364_),
    .Y(net218));
 sky130_fd_sc_hd__nor2_1 _1926_ (.A(_0322_),
    .B(_0256_),
    .Y(_0365_));
 sky130_fd_sc_hd__a31oi_2 _1927_ (.A1(_0267_),
    .A2(_0321_),
    .A3(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[28] ),
    .B1(_0365_),
    .Y(_0366_));
 sky130_fd_sc_hd__nand2_1 _1928_ (.A(_0336_),
    .B(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[28] ),
    .Y(_0367_));
 sky130_fd_sc_hd__o21ai_2 _1929_ (.A1(_0351_),
    .A2(_0366_),
    .B1(_0367_),
    .Y(net219));
 sky130_fd_sc_hd__mux2i_2 _1930_ (.A0(_0260_),
    .A1(_0133_),
    .S(_0321_),
    .Y(_0368_));
 sky130_fd_sc_hd__nand2_1 _1931_ (.A(_0336_),
    .B(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[29] ),
    .Y(_0369_));
 sky130_fd_sc_hd__o21ai_2 _1932_ (.A1(_0351_),
    .A2(_0368_),
    .B1(_0369_),
    .Y(net220));
 sky130_fd_sc_hd__mux2_1 _1933_ (.A0(_0873_),
    .A1(_0874_),
    .S(_0773_),
    .X(_0370_));
 sky130_fd_sc_hd__nand2_1 _1934_ (.A(_0336_),
    .B(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[2] ),
    .Y(_0371_));
 sky130_fd_sc_hd__o21ai_4 _1935_ (.A1(_0351_),
    .A2(_0370_),
    .B1(_0371_),
    .Y(net221));
 sky130_fd_sc_hd__nor2_1 _1936_ (.A(_0772_),
    .B(_0143_),
    .Y(_0372_));
 sky130_fd_sc_hd__a21oi_1 _1937_ (.A1(_0304_),
    .A2(_0142_),
    .B1(_0372_),
    .Y(_0373_));
 sky130_fd_sc_hd__nand2_1 _1938_ (.A(_0303_),
    .B(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[30] ),
    .Y(_0374_));
 sky130_fd_sc_hd__o21ai_2 _1939_ (.A1(_0351_),
    .A2(_0373_),
    .B1(_0374_),
    .Y(net222));
 sky130_fd_sc_hd__nand2_1 _1940_ (.A(_0305_),
    .B(_0153_),
    .Y(_0375_));
 sky130_fd_sc_hd__o21ai_1 _1941_ (.A1(_0304_),
    .A2(_0149_),
    .B1(_0375_),
    .Y(_0376_));
 sky130_fd_sc_hd__nand2_1 _1942_ (.A(_0303_),
    .B(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[31] ),
    .Y(_0377_));
 sky130_fd_sc_hd__o21ai_4 _1943_ (.A1(_0351_),
    .A2(_0376_),
    .B1(_0377_),
    .Y(net223));
 sky130_fd_sc_hd__o211ai_1 _1944_ (.A1(_0858_),
    .A2(_0868_),
    .B1(_0856_),
    .C1(_0305_),
    .Y(_0378_));
 sky130_fd_sc_hd__o21ai_1 _1945_ (.A1(_0304_),
    .A2(_0862_),
    .B1(_0378_),
    .Y(_0379_));
 sky130_fd_sc_hd__nand2_1 _1946_ (.A(_0303_),
    .B(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[3] ),
    .Y(_0380_));
 sky130_fd_sc_hd__o21ai_4 _1947_ (.A1(_0351_),
    .A2(_0379_),
    .B1(_0380_),
    .Y(net224));
 sky130_fd_sc_hd__nor2_1 _1948_ (.A(_0305_),
    .B(_0944_),
    .Y(_0381_));
 sky130_fd_sc_hd__a211oi_4 _1949_ (.A1(net149),
    .A2(_0867_),
    .B1(_0940_),
    .C1(_0321_),
    .Y(_0382_));
 sky130_fd_sc_hd__nand2_1 _1950_ (.A(_0309_),
    .B(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[4] ),
    .Y(_0383_));
 sky130_fd_sc_hd__o31ai_4 _1951_ (.A1(_0308_),
    .A2(_0381_),
    .A3(_0382_),
    .B1(_0383_),
    .Y(net225));
 sky130_fd_sc_hd__a21oi_1 _1952_ (.A1(net150),
    .A2(_0867_),
    .B1(_0957_),
    .Y(_0384_));
 sky130_fd_sc_hd__nand2_1 _1953_ (.A(_0322_),
    .B(_0953_),
    .Y(_0385_));
 sky130_fd_sc_hd__o21ai_1 _1954_ (.A1(_0322_),
    .A2(_0384_),
    .B1(_0385_),
    .Y(_0386_));
 sky130_fd_sc_hd__mux2_2 _1955_ (.A0(_0386_),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[5] ),
    .S(_0308_),
    .X(net226));
 sky130_fd_sc_hd__a21oi_1 _1956_ (.A1(net151),
    .A2(_0867_),
    .B1(_0951_),
    .Y(_0387_));
 sky130_fd_sc_hd__nand2_1 _1957_ (.A(_0322_),
    .B(_0947_),
    .Y(_0388_));
 sky130_fd_sc_hd__o21ai_0 _1958_ (.A1(_0322_),
    .A2(_0387_),
    .B1(_0388_),
    .Y(_0389_));
 sky130_fd_sc_hd__mux2_2 _1959_ (.A0(_0389_),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[6] ),
    .S(_0308_),
    .X(net227));
 sky130_fd_sc_hd__a2111oi_4 _1960_ (.A1(_0932_),
    .A2(_0933_),
    .B1(_0934_),
    .C1(_0935_),
    .D1(_0322_),
    .Y(_0390_));
 sky130_fd_sc_hd__a21oi_2 _1961_ (.A1(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[7] ),
    .A2(_0327_),
    .B1(_0390_),
    .Y(_0391_));
 sky130_fd_sc_hd__nand2_1 _1962_ (.A(_0303_),
    .B(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[7] ),
    .Y(_0392_));
 sky130_fd_sc_hd__o21ai_4 _1963_ (.A1(_0351_),
    .A2(_0391_),
    .B1(_0392_),
    .Y(net228));
 sky130_fd_sc_hd__a22oi_4 _1964_ (.A1(_0305_),
    .A2(_0164_),
    .B1(_0327_),
    .B2(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[8] ),
    .Y(_0393_));
 sky130_fd_sc_hd__nand2_1 _1965_ (.A(_0303_),
    .B(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[8] ),
    .Y(_0394_));
 sky130_fd_sc_hd__o21ai_4 _1966_ (.A1(_0308_),
    .A2(_0393_),
    .B1(_0394_),
    .Y(net229));
 sky130_fd_sc_hd__nor2_1 _1967_ (.A(net29),
    .B(_0912_),
    .Y(_0395_));
 sky130_fd_sc_hd__nor2_1 _1968_ (.A(_0395_),
    .B(_0965_),
    .Y(_0396_));
 sky130_fd_sc_hd__nor2_1 _1969_ (.A(_0772_),
    .B(_0967_),
    .Y(_0397_));
 sky130_fd_sc_hd__a21oi_2 _1970_ (.A1(_0304_),
    .A2(_0396_),
    .B1(_0397_),
    .Y(_0398_));
 sky130_fd_sc_hd__nand2_1 _1971_ (.A(_0303_),
    .B(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[9] ),
    .Y(_0399_));
 sky130_fd_sc_hd__o21ai_4 _1972_ (.A1(_0308_),
    .A2(_0398_),
    .B1(_0399_),
    .Y(net230));
 sky130_fd_sc_hd__nor2_1 _1973_ (.A(_0778_),
    .B(_0838_),
    .Y(_0400_));
 sky130_fd_sc_hd__a221o_1 _1974_ (.A1(_0893_),
    .A2(_0838_),
    .B1(_0892_),
    .B2(net315),
    .C1(_0400_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[0] ));
 sky130_fd_sc_hd__a31oi_1 _1975_ (.A1(_0893_),
    .A2(net315),
    .A3(_0892_),
    .B1(\gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1] ),
    .Y(_0401_));
 sky130_fd_sc_hd__nor2_1 _1976_ (.A(_0894_),
    .B(_0401_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[1] ));
 sky130_fd_sc_hd__nand2_1 _1977_ (.A(net157),
    .B(net315),
    .Y(_0402_));
 sky130_fd_sc_hd__nand2_1 _1978_ (.A(_0893_),
    .B(net190),
    .Y(_0403_));
 sky130_fd_sc_hd__o21ai_0 _1979_ (.A1(_0893_),
    .A2(_0402_),
    .B1(_0403_),
    .Y(_0404_));
 sky130_fd_sc_hd__nor2b_1 _1980_ (.A(\gen_prefetch_buffer.prefetch_buffer_i.rdata_pmp_err_q[1] ),
    .B_N(_0893_),
    .Y(_0405_));
 sky130_fd_sc_hd__o21ai_0 _1981_ (.A1(\gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1] ),
    .A2(_0402_),
    .B1(_0405_),
    .Y(_0406_));
 sky130_fd_sc_hd__o21a_1 _1982_ (.A1(\gen_prefetch_buffer.prefetch_buffer_i.rdata_pmp_err_q[0] ),
    .A2(_0404_),
    .B1(_0406_),
    .X(\gen_prefetch_buffer.prefetch_buffer_i.rdata_pmp_err_s[0] ));
 sky130_fd_sc_hd__a41oi_1 _1983_ (.A1(_0893_),
    .A2(_0778_),
    .A3(net157),
    .A4(net315),
    .B1(\gen_prefetch_buffer.prefetch_buffer_i.rdata_pmp_err_q[1] ),
    .Y(_0407_));
 sky130_fd_sc_hd__nor2_1 _1984_ (.A(_0894_),
    .B(_0407_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.rdata_pmp_err_s[1] ));
 sky130_fd_sc_hd__nor2_8 _1985_ (.A(_0864_),
    .B(_0892_),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ));
 sky130_fd_sc_hd__nor2b_1 _1986_ (.A(_0892_),
    .B_N(net315),
    .Y(\gen_prefetch_buffer.prefetch_buffer_i.valid_req_d ));
 sky130_fd_sc_hd__or3_2 _1987_ (.A(_0893_),
    .B(\gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1] ),
    .C(net315),
    .X(net199));
 sky130_fd_sc_hd__buf_8 _1988_ (.A(_0752_),
    .X(_0408_));
 sky130_fd_sc_hd__buf_4 _1989_ (.A(_0408_),
    .X(_0409_));
 sky130_fd_sc_hd__buf_4 _1990_ (.A(_0758_),
    .X(_0410_));
 sky130_fd_sc_hd__buf_4 _1991_ (.A(_0795_),
    .X(_0411_));
 sky130_fd_sc_hd__buf_4 _1992_ (.A(_0806_),
    .X(_0412_));
 sky130_fd_sc_hd__nor2_1 _1993_ (.A(_0802_),
    .B(_0803_),
    .Y(_0413_));
 sky130_fd_sc_hd__nor4b_4 _1994_ (.A(_0811_),
    .B(\compressed_decoder_i.instr_i[3] ),
    .C(\compressed_decoder_i.instr_i[4] ),
    .D_N(_0413_),
    .Y(_0414_));
 sky130_fd_sc_hd__buf_2 _1995_ (.A(_0414_),
    .X(_0415_));
 sky130_fd_sc_hd__nand2_8 _1996_ (.A(_0788_),
    .B(_0833_),
    .Y(_0416_));
 sky130_fd_sc_hd__a31oi_1 _1997_ (.A1(_0411_),
    .A2(_0412_),
    .A3(_0415_),
    .B1(_0416_),
    .Y(_0417_));
 sky130_fd_sc_hd__buf_6 _1998_ (.A(_0831_),
    .X(_0418_));
 sky130_fd_sc_hd__nand2_1 _1999_ (.A(_0411_),
    .B(_0418_),
    .Y(_0419_));
 sky130_fd_sc_hd__nor4_4 _2000_ (.A(_0800_),
    .B(_0801_),
    .C(_0813_),
    .D(\compressed_decoder_i.instr_i[9] ),
    .Y(_0420_));
 sky130_fd_sc_hd__and2_2 _2001_ (.A(_0816_),
    .B(_0420_),
    .X(_0421_));
 sky130_fd_sc_hd__nor2_1 _2002_ (.A(_0412_),
    .B(_0419_),
    .Y(_0422_));
 sky130_fd_sc_hd__a211oi_1 _2003_ (.A1(_0419_),
    .A2(_0421_),
    .B1(_0422_),
    .C1(\compressed_decoder_i.instr_i[13] ),
    .Y(_0423_));
 sky130_fd_sc_hd__clkinv_2 _2004_ (.A(\compressed_decoder_i.instr_i[11] ),
    .Y(_0424_));
 sky130_fd_sc_hd__nor3b_1 _2005_ (.A(_0790_),
    .B(_0796_),
    .C_N(_0832_),
    .Y(_0425_));
 sky130_fd_sc_hd__buf_4 _2006_ (.A(_0425_),
    .X(_0426_));
 sky130_fd_sc_hd__o211ai_1 _2007_ (.A1(_0424_),
    .A2(_0801_),
    .B1(\compressed_decoder_i.instr_i[12] ),
    .C1(_0426_),
    .Y(_0427_));
 sky130_fd_sc_hd__nand2_1 _2008_ (.A(_0790_),
    .B(_0797_),
    .Y(_0428_));
 sky130_fd_sc_hd__nor2_2 _2009_ (.A(_0833_),
    .B(_0428_),
    .Y(_0429_));
 sky130_fd_sc_hd__nand3_1 _2010_ (.A(_0806_),
    .B(_0415_),
    .C(_0429_),
    .Y(_0430_));
 sky130_fd_sc_hd__nand2_8 _2011_ (.A(_0788_),
    .B(_0418_),
    .Y(_0431_));
 sky130_fd_sc_hd__nor2_8 _2012_ (.A(_0797_),
    .B(_0431_),
    .Y(_0432_));
 sky130_fd_sc_hd__nor3_4 _2013_ (.A(_0802_),
    .B(_0803_),
    .C(_0807_),
    .Y(_0433_));
 sky130_fd_sc_hd__nand2b_4 _2014_ (.A_N(_0796_),
    .B(_0832_),
    .Y(_0434_));
 sky130_fd_sc_hd__nand2_8 _2015_ (.A(_0788_),
    .B(_0434_),
    .Y(_0435_));
 sky130_fd_sc_hd__a311oi_4 _2016_ (.A1(_0421_),
    .A2(_0432_),
    .A3(_0433_),
    .B1(_0435_),
    .C1(_0758_),
    .Y(_0436_));
 sky130_fd_sc_hd__a311o_1 _2017_ (.A1(_0410_),
    .A2(_0427_),
    .A3(_0430_),
    .B1(_0436_),
    .C1(\compressed_decoder_i.instr_i[1] ),
    .X(_0437_));
 sky130_fd_sc_hd__o41ai_1 _2018_ (.A1(_0409_),
    .A2(_0410_),
    .A3(_0417_),
    .A4(_0423_),
    .B1(_0437_),
    .Y(\compressed_decoder_i.illegal_instr_o ));
 sky130_fd_sc_hd__nor2_2 _2019_ (.A(_0753_),
    .B(_0434_),
    .Y(_0438_));
 sky130_fd_sc_hd__o21ai_2 _2020_ (.A1(_0790_),
    .A2(_0438_),
    .B1(_0757_),
    .Y(\compressed_decoder_i.instr_o[0] ));
 sky130_fd_sc_hd__nand2_1 _2021_ (.A(_0415_),
    .B(_0426_),
    .Y(_0439_));
 sky130_fd_sc_hd__nor3_1 _2022_ (.A(_0409_),
    .B(_0410_),
    .C(_0439_),
    .Y(_0440_));
 sky130_fd_sc_hd__nand2_4 _2023_ (.A(_0790_),
    .B(_0795_),
    .Y(_0441_));
 sky130_fd_sc_hd__nand2_8 _2024_ (.A(_0408_),
    .B(_0758_),
    .Y(_0442_));
 sky130_fd_sc_hd__o21ai_0 _2025_ (.A1(_0441_),
    .A2(_0442_),
    .B1(\compressed_decoder_i.instr_i[10] ),
    .Y(_0443_));
 sky130_fd_sc_hd__buf_4 _2026_ (.A(_0418_),
    .X(_0444_));
 sky130_fd_sc_hd__nand2_1 _2027_ (.A(_0410_),
    .B(_0434_),
    .Y(_0445_));
 sky130_fd_sc_hd__buf_4 _2028_ (.A(_0788_),
    .X(_0446_));
 sky130_fd_sc_hd__buf_6 _2029_ (.A(_0446_),
    .X(_0447_));
 sky130_fd_sc_hd__o2111ai_1 _2030_ (.A1(_0410_),
    .A2(_0444_),
    .B1(_0445_),
    .C1(_0447_),
    .D1(_0409_),
    .Y(_0448_));
 sky130_fd_sc_hd__o21ai_1 _2031_ (.A1(_0440_),
    .A2(_0443_),
    .B1(_0448_),
    .Y(\compressed_decoder_i.instr_o[10] ));
 sky130_fd_sc_hd__nand2_1 _2032_ (.A(\compressed_decoder_i.instr_i[1] ),
    .B(_0439_),
    .Y(_0449_));
 sky130_fd_sc_hd__nand2_1 _2033_ (.A(\compressed_decoder_i.instr_i[10] ),
    .B(_0808_),
    .Y(_0450_));
 sky130_fd_sc_hd__a21oi_1 _2034_ (.A1(\compressed_decoder_i.instr_i[15] ),
    .A2(_0450_),
    .B1(\compressed_decoder_i.instr_i[13] ),
    .Y(_0451_));
 sky130_fd_sc_hd__nor2_8 _2035_ (.A(_0790_),
    .B(_0832_),
    .Y(_0452_));
 sky130_fd_sc_hd__nor2_1 _2036_ (.A(_0754_),
    .B(_0452_),
    .Y(_0453_));
 sky130_fd_sc_hd__o32ai_1 _2037_ (.A1(\compressed_decoder_i.instr_i[14] ),
    .A2(_0442_),
    .A3(_0451_),
    .B1(_0453_),
    .B2(\compressed_decoder_i.instr_i[0] ),
    .Y(_0454_));
 sky130_fd_sc_hd__a21oi_1 _2038_ (.A1(_0449_),
    .A2(_0454_),
    .B1(_0424_),
    .Y(\compressed_decoder_i.instr_o[11] ));
 sky130_fd_sc_hd__nand2_8 _2039_ (.A(_0795_),
    .B(_0452_),
    .Y(_0455_));
 sky130_fd_sc_hd__nor2_1 _2040_ (.A(_0753_),
    .B(_0757_),
    .Y(_0456_));
 sky130_fd_sc_hd__buf_6 _2041_ (.A(_0456_),
    .X(_0457_));
 sky130_fd_sc_hd__nand2_4 _2042_ (.A(_0455_),
    .B(_0457_),
    .Y(_0458_));
 sky130_fd_sc_hd__nor2_4 _2043_ (.A(_0797_),
    .B(_0418_),
    .Y(_0459_));
 sky130_fd_sc_hd__nand2_8 _2044_ (.A(\compressed_decoder_i.instr_i[11] ),
    .B(_0801_),
    .Y(_0460_));
 sky130_fd_sc_hd__a21oi_1 _2045_ (.A1(\compressed_decoder_i.instr_i[5] ),
    .A2(\compressed_decoder_i.instr_i[6] ),
    .B1(_0460_),
    .Y(_0461_));
 sky130_fd_sc_hd__o21ai_0 _2046_ (.A1(_0791_),
    .A2(_0461_),
    .B1(_0412_),
    .Y(_0462_));
 sky130_fd_sc_hd__nand2_4 _2047_ (.A(\compressed_decoder_i.instr_i[8] ),
    .B(_0420_),
    .Y(_0463_));
 sky130_fd_sc_hd__nand2_1 _2048_ (.A(_0798_),
    .B(_0418_),
    .Y(_0464_));
 sky130_fd_sc_hd__a21oi_1 _2049_ (.A1(\compressed_decoder_i.instr_i[2] ),
    .A2(_0463_),
    .B1(_0464_),
    .Y(_0465_));
 sky130_fd_sc_hd__a211oi_1 _2050_ (.A1(_0411_),
    .A2(_0412_),
    .B1(_0465_),
    .C1(_0447_),
    .Y(_0466_));
 sky130_fd_sc_hd__a21oi_1 _2051_ (.A1(_0459_),
    .A2(_0462_),
    .B1(_0466_),
    .Y(_0467_));
 sky130_fd_sc_hd__buf_4 _2052_ (.A(_0757_),
    .X(_0468_));
 sky130_fd_sc_hd__nand2_2 _2053_ (.A(_0757_),
    .B(_0446_),
    .Y(_0469_));
 sky130_fd_sc_hd__o22ai_1 _2054_ (.A1(_0468_),
    .A2(_0412_),
    .B1(_0419_),
    .B2(_0469_),
    .Y(_0470_));
 sky130_fd_sc_hd__nand2_1 _2055_ (.A(\compressed_decoder_i.instr_i[1] ),
    .B(_0470_),
    .Y(_0471_));
 sky130_fd_sc_hd__o211ai_1 _2056_ (.A1(\compressed_decoder_i.instr_i[13] ),
    .A2(_0438_),
    .B1(\compressed_decoder_i.instr_i[12] ),
    .C1(_0468_),
    .Y(_0472_));
 sky130_fd_sc_hd__o211ai_1 _2057_ (.A1(_0458_),
    .A2(_0467_),
    .B1(_0471_),
    .C1(_0472_),
    .Y(\compressed_decoder_i.instr_o[12] ));
 sky130_fd_sc_hd__nor2_2 _2058_ (.A(_0790_),
    .B(_0798_),
    .Y(_0473_));
 sky130_fd_sc_hd__nor2_4 _2059_ (.A(_0432_),
    .B(_0442_),
    .Y(_0474_));
 sky130_fd_sc_hd__clkinv_2 _2060_ (.A(\compressed_decoder_i.instr_i[3] ),
    .Y(_0475_));
 sky130_fd_sc_hd__nand2_2 _2061_ (.A(_0429_),
    .B(_0463_),
    .Y(_0476_));
 sky130_fd_sc_hd__clkinvlp_4 _2062_ (.A(\compressed_decoder_i.instr_i[6] ),
    .Y(_0477_));
 sky130_fd_sc_hd__o21ai_0 _2063_ (.A1(_0477_),
    .A2(_0808_),
    .B1(_0801_),
    .Y(_0478_));
 sky130_fd_sc_hd__a32oi_1 _2064_ (.A1(\compressed_decoder_i.instr_i[11] ),
    .A2(_0426_),
    .A3(_0478_),
    .B1(\compressed_decoder_i.instr_i[12] ),
    .B2(_0791_),
    .Y(_0479_));
 sky130_fd_sc_hd__o22ai_1 _2065_ (.A1(_0475_),
    .A2(_0476_),
    .B1(_0479_),
    .B2(\compressed_decoder_i.instr_i[14] ),
    .Y(_0480_));
 sky130_fd_sc_hd__nand2_1 _2066_ (.A(_0474_),
    .B(_0480_),
    .Y(_0481_));
 sky130_fd_sc_hd__o221ai_2 _2067_ (.A1(_0409_),
    .A2(_0447_),
    .B1(_0473_),
    .B2(\compressed_decoder_i.instr_i[0] ),
    .C1(_0481_),
    .Y(\compressed_decoder_i.instr_o[13] ));
 sky130_fd_sc_hd__nand3_1 _2068_ (.A(\compressed_decoder_i.instr_i[4] ),
    .B(_0429_),
    .C(_0463_),
    .Y(_0482_));
 sky130_fd_sc_hd__nor2_1 _2069_ (.A(\compressed_decoder_i.instr_i[12] ),
    .B(_0413_),
    .Y(_0483_));
 sky130_fd_sc_hd__o21ai_0 _2070_ (.A1(_0460_),
    .A2(_0483_),
    .B1(_0426_),
    .Y(_0484_));
 sky130_fd_sc_hd__nor2_2 _2071_ (.A(_0446_),
    .B(_0798_),
    .Y(_0485_));
 sky130_fd_sc_hd__a21oi_1 _2072_ (.A1(\compressed_decoder_i.instr_i[12] ),
    .A2(_0485_),
    .B1(_0442_),
    .Y(_0486_));
 sky130_fd_sc_hd__o21ai_0 _2073_ (.A1(\compressed_decoder_i.instr_i[14] ),
    .A2(_0453_),
    .B1(\compressed_decoder_i.instr_i[0] ),
    .Y(_0487_));
 sky130_fd_sc_hd__a32oi_2 _2074_ (.A1(_0482_),
    .A2(_0484_),
    .A3(_0486_),
    .B1(_0487_),
    .B2(_0428_),
    .Y(\compressed_decoder_i.instr_o[14] ));
 sky130_fd_sc_hd__nor2b_4 _2075_ (.A(_0790_),
    .B_N(_0797_),
    .Y(_0488_));
 sky130_fd_sc_hd__nand2_1 _2076_ (.A(\compressed_decoder_i.instr_i[7] ),
    .B(_0488_),
    .Y(_0489_));
 sky130_fd_sc_hd__o21ai_0 _2077_ (.A1(_0444_),
    .A2(_0488_),
    .B1(_0489_),
    .Y(_0490_));
 sky130_fd_sc_hd__o31ai_4 _2078_ (.A1(_0808_),
    .A2(_0418_),
    .A3(_0414_),
    .B1(_0473_),
    .Y(_0491_));
 sky130_fd_sc_hd__inv_1 _2079_ (.A(_0813_),
    .Y(_0492_));
 sky130_fd_sc_hd__o221ai_1 _2080_ (.A1(_0447_),
    .A2(_0444_),
    .B1(_0491_),
    .B2(_0492_),
    .C1(\compressed_decoder_i.instr_i[1] ),
    .Y(_0493_));
 sky130_fd_sc_hd__o21ai_0 _2081_ (.A1(\compressed_decoder_i.instr_i[1] ),
    .A2(_0490_),
    .B1(_0493_),
    .Y(_0494_));
 sky130_fd_sc_hd__a21oi_1 _2082_ (.A1(_0446_),
    .A2(_0460_),
    .B1(_0806_),
    .Y(_0495_));
 sky130_fd_sc_hd__o21ai_0 _2083_ (.A1(_0452_),
    .A2(_0495_),
    .B1(_0411_),
    .Y(_0496_));
 sky130_fd_sc_hd__nand3_1 _2084_ (.A(_0802_),
    .B(_0429_),
    .C(_0463_),
    .Y(_0497_));
 sky130_fd_sc_hd__a221oi_1 _2085_ (.A1(_0492_),
    .A2(_0432_),
    .B1(_0496_),
    .B2(_0497_),
    .C1(_0754_),
    .Y(_0498_));
 sky130_fd_sc_hd__nand2_2 _2086_ (.A(_0797_),
    .B(_0833_),
    .Y(_0499_));
 sky130_fd_sc_hd__a21oi_1 _2087_ (.A1(_0802_),
    .A2(\compressed_decoder_i.instr_i[6] ),
    .B1(_0807_),
    .Y(_0500_));
 sky130_fd_sc_hd__o21ai_2 _2088_ (.A1(_0460_),
    .A2(_0500_),
    .B1(_0425_),
    .Y(_0501_));
 sky130_fd_sc_hd__nand2_1 _2089_ (.A(_0499_),
    .B(_0501_),
    .Y(_0502_));
 sky130_fd_sc_hd__nand3_2 _2090_ (.A(_0802_),
    .B(\compressed_decoder_i.instr_i[6] ),
    .C(_0806_),
    .Y(_0503_));
 sky130_fd_sc_hd__nor2_1 _2091_ (.A(_0416_),
    .B(_0503_),
    .Y(_0504_));
 sky130_fd_sc_hd__o211a_1 _2092_ (.A1(_0502_),
    .A2(_0504_),
    .B1(_0408_),
    .C1(\compressed_decoder_i.instr_i[7] ),
    .X(_0505_));
 sky130_fd_sc_hd__a2111oi_0 _2093_ (.A1(_0754_),
    .A2(\compressed_decoder_i.instr_i[15] ),
    .B1(_0498_),
    .C1(_0505_),
    .D1(_0468_),
    .Y(_0506_));
 sky130_fd_sc_hd__a21oi_1 _2094_ (.A1(_0468_),
    .A2(_0494_),
    .B1(_0506_),
    .Y(\compressed_decoder_i.instr_o[15] ));
 sky130_fd_sc_hd__nand2_1 _2095_ (.A(_0836_),
    .B(_0292_),
    .Y(_0507_));
 sky130_fd_sc_hd__o21ai_4 _2096_ (.A1(_0836_),
    .A2(_0755_),
    .B1(_0507_),
    .Y(_0508_));
 sky130_fd_sc_hd__nand2_4 _2097_ (.A(_0753_),
    .B(_0758_),
    .Y(\compressed_decoder_i.is_compressed_o ));
 sky130_fd_sc_hd__nor2_1 _2098_ (.A(_0508_),
    .B(\compressed_decoder_i.is_compressed_o ),
    .Y(_0509_));
 sky130_fd_sc_hd__nand2_4 _2099_ (.A(_0408_),
    .B(_0757_),
    .Y(_0510_));
 sky130_fd_sc_hd__a221oi_1 _2100_ (.A1(_0816_),
    .A2(_0488_),
    .B1(_0435_),
    .B2(_0508_),
    .C1(_0510_),
    .Y(_0511_));
 sky130_fd_sc_hd__or3b_4 _2101_ (.A(_0789_),
    .B(_0796_),
    .C_N(_0832_),
    .X(_0512_));
 sky130_fd_sc_hd__nor3_1 _2102_ (.A(\compressed_decoder_i.instr_i[12] ),
    .B(_0415_),
    .C(_0512_),
    .Y(_0513_));
 sky130_fd_sc_hd__nand2_4 _2103_ (.A(_0753_),
    .B(_0757_),
    .Y(_0514_));
 sky130_fd_sc_hd__a21o_1 _2104_ (.A1(_0791_),
    .A2(_0508_),
    .B1(_0514_),
    .X(_0515_));
 sky130_fd_sc_hd__a211oi_1 _2105_ (.A1(_0816_),
    .A2(_0473_),
    .B1(_0513_),
    .C1(_0515_),
    .Y(_0516_));
 sky130_fd_sc_hd__nor3_1 _2106_ (.A(_0509_),
    .B(_0511_),
    .C(_0516_),
    .Y(_0517_));
 sky130_fd_sc_hd__nor2_2 _2107_ (.A(_0433_),
    .B(_0512_),
    .Y(_0518_));
 sky130_fd_sc_hd__nand3_4 _2108_ (.A(\compressed_decoder_i.instr_i[11] ),
    .B(_0801_),
    .C(_0807_),
    .Y(_0519_));
 sky130_fd_sc_hd__o22ai_1 _2109_ (.A1(_0816_),
    .A2(_0503_),
    .B1(_0508_),
    .B2(_0519_),
    .Y(_0520_));
 sky130_fd_sc_hd__nand2_1 _2110_ (.A(_0797_),
    .B(\compressed_decoder_i.instr_i[6] ),
    .Y(_0521_));
 sky130_fd_sc_hd__o22ai_1 _2111_ (.A1(_0797_),
    .A2(_0806_),
    .B1(_0833_),
    .B2(_0521_),
    .Y(_0522_));
 sky130_fd_sc_hd__a221o_1 _2112_ (.A1(_0518_),
    .A2(_0520_),
    .B1(_0522_),
    .B2(_0790_),
    .C1(_0432_),
    .X(_0523_));
 sky130_fd_sc_hd__nand2_1 _2113_ (.A(_0474_),
    .B(_0523_),
    .Y(_0524_));
 sky130_fd_sc_hd__nor3_4 _2114_ (.A(_0446_),
    .B(_0464_),
    .C(_0463_),
    .Y(_0525_));
 sky130_fd_sc_hd__o311ai_1 _2115_ (.A1(_0502_),
    .A2(_0523_),
    .A3(_0525_),
    .B1(_0457_),
    .C1(\compressed_decoder_i.instr_i[8] ),
    .Y(_0526_));
 sky130_fd_sc_hd__nand3_1 _2116_ (.A(_0517_),
    .B(_0524_),
    .C(_0526_),
    .Y(\compressed_decoder_i.instr_o[16] ));
 sky130_fd_sc_hd__mux2i_4 _2117_ (.A0(_0748_),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[1] ),
    .S(_0836_),
    .Y(_0527_));
 sky130_fd_sc_hd__nor2_4 _2118_ (.A(_0408_),
    .B(_0758_),
    .Y(_0528_));
 sky130_fd_sc_hd__o22ai_1 _2119_ (.A1(_0820_),
    .A2(_0491_),
    .B1(_0527_),
    .B2(_0447_),
    .Y(_0529_));
 sky130_fd_sc_hd__nand2_1 _2120_ (.A(_0528_),
    .B(_0529_),
    .Y(_0530_));
 sky130_fd_sc_hd__nor2_2 _2121_ (.A(_0753_),
    .B(_0758_),
    .Y(_0531_));
 sky130_fd_sc_hd__nand2_4 _2122_ (.A(_0446_),
    .B(_0798_),
    .Y(_0532_));
 sky130_fd_sc_hd__nor2_2 _2123_ (.A(_0791_),
    .B(_0459_),
    .Y(_0533_));
 sky130_fd_sc_hd__o22ai_1 _2124_ (.A1(_0820_),
    .A2(_0532_),
    .B1(_0533_),
    .B2(_0527_),
    .Y(_0534_));
 sky130_fd_sc_hd__nand2_1 _2125_ (.A(_0531_),
    .B(_0534_),
    .Y(_0535_));
 sky130_fd_sc_hd__o22ai_1 _2126_ (.A1(_0820_),
    .A2(_0503_),
    .B1(_0519_),
    .B2(_0527_),
    .Y(_0536_));
 sky130_fd_sc_hd__nand2_1 _2127_ (.A(_0790_),
    .B(_0807_),
    .Y(_0537_));
 sky130_fd_sc_hd__and2_4 _2128_ (.A(_0796_),
    .B(_0832_),
    .X(_0538_));
 sky130_fd_sc_hd__a311o_1 _2129_ (.A1(_0797_),
    .A2(\compressed_decoder_i.instr_i[8] ),
    .A3(_0420_),
    .B1(_0537_),
    .C1(_0538_),
    .X(_0539_));
 sky130_fd_sc_hd__nand2_2 _2130_ (.A(_0455_),
    .B(_0539_),
    .Y(_0540_));
 sky130_fd_sc_hd__a221o_1 _2131_ (.A1(\compressed_decoder_i.instr_i[9] ),
    .A2(_0502_),
    .B1(_0518_),
    .B2(_0536_),
    .C1(_0540_),
    .X(_0541_));
 sky130_fd_sc_hd__nand2_1 _2132_ (.A(_0820_),
    .B(_0432_),
    .Y(_0542_));
 sky130_fd_sc_hd__nand3_1 _2133_ (.A(_0457_),
    .B(_0541_),
    .C(_0542_),
    .Y(_0543_));
 sky130_fd_sc_hd__o2111ai_1 _2134_ (.A1(\compressed_decoder_i.is_compressed_o ),
    .A2(_0527_),
    .B1(_0530_),
    .C1(_0535_),
    .D1(_0543_),
    .Y(\compressed_decoder_i.instr_o[17] ));
 sky130_fd_sc_hd__nor2_4 _2135_ (.A(_0806_),
    .B(_0460_),
    .Y(_0544_));
 sky130_fd_sc_hd__nand2_1 _2136_ (.A(_0751_),
    .B(_0809_),
    .Y(_0545_));
 sky130_fd_sc_hd__o21ai_4 _2137_ (.A1(_0751_),
    .A2(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[2] ),
    .B1(_0545_),
    .Y(_0546_));
 sky130_fd_sc_hd__a21oi_1 _2138_ (.A1(_0544_),
    .A2(_0546_),
    .B1(_0416_),
    .Y(_0547_));
 sky130_fd_sc_hd__inv_1 _2139_ (.A(_0801_),
    .Y(_0548_));
 sky130_fd_sc_hd__nand2_1 _2140_ (.A(_0548_),
    .B(_0432_),
    .Y(_0549_));
 sky130_fd_sc_hd__o311a_1 _2141_ (.A1(_0538_),
    .A2(_0540_),
    .A3(_0547_),
    .B1(_0549_),
    .C1(_0457_),
    .X(_0550_));
 sky130_fd_sc_hd__nand2_2 _2142_ (.A(_0754_),
    .B(_0469_),
    .Y(_0551_));
 sky130_fd_sc_hd__nand2_1 _2143_ (.A(_0468_),
    .B(\compressed_decoder_i.instr_i[10] ),
    .Y(_0552_));
 sky130_fd_sc_hd__o221ai_1 _2144_ (.A1(_0546_),
    .A2(_0551_),
    .B1(_0552_),
    .B2(_0491_),
    .C1(_0510_),
    .Y(_0553_));
 sky130_fd_sc_hd__nor2_2 _2145_ (.A(_0488_),
    .B(_0510_),
    .Y(_0554_));
 sky130_fd_sc_hd__o21ai_0 _2146_ (.A1(_0452_),
    .A2(_0546_),
    .B1(_0554_),
    .Y(_0555_));
 sky130_fd_sc_hd__o21a_1 _2147_ (.A1(_0550_),
    .A2(_0553_),
    .B1(_0555_),
    .X(\compressed_decoder_i.instr_o[18] ));
 sky130_fd_sc_hd__mux2_1 _2148_ (.A0(net168),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[19] ),
    .S(_0877_),
    .X(_0556_));
 sky130_fd_sc_hd__nand2_1 _2149_ (.A(_0887_),
    .B(_0822_),
    .Y(_0557_));
 sky130_fd_sc_hd__o21ai_4 _2150_ (.A1(_0887_),
    .A2(_0556_),
    .B1(_0557_),
    .Y(_0558_));
 sky130_fd_sc_hd__o22ai_1 _2151_ (.A1(_0424_),
    .A2(_0491_),
    .B1(_0558_),
    .B2(_0447_),
    .Y(_0559_));
 sky130_fd_sc_hd__nand2_1 _2152_ (.A(_0528_),
    .B(_0559_),
    .Y(_0560_));
 sky130_fd_sc_hd__o211ai_1 _2153_ (.A1(\compressed_decoder_i.instr_i[11] ),
    .A2(_0455_),
    .B1(_0457_),
    .C1(_0540_),
    .Y(_0561_));
 sky130_fd_sc_hd__a21oi_1 _2154_ (.A1(_0408_),
    .A2(_0435_),
    .B1(_0758_),
    .Y(_0562_));
 sky130_fd_sc_hd__a21oi_1 _2155_ (.A1(_0426_),
    .A2(_0544_),
    .B1(_0442_),
    .Y(_0563_));
 sky130_fd_sc_hd__nor2_2 _2156_ (.A(_0562_),
    .B(_0563_),
    .Y(_0564_));
 sky130_fd_sc_hd__nand2b_1 _2157_ (.A_N(_0558_),
    .B(_0564_),
    .Y(_0565_));
 sky130_fd_sc_hd__nand3_1 _2158_ (.A(_0560_),
    .B(_0561_),
    .C(_0565_),
    .Y(\compressed_decoder_i.instr_o[19] ));
 sky130_fd_sc_hd__o21ai_0 _2159_ (.A1(\compressed_decoder_i.instr_i[13] ),
    .A2(_0519_),
    .B1(\compressed_decoder_i.instr_i[0] ),
    .Y(_0566_));
 sky130_fd_sc_hd__nand3_1 _2160_ (.A(_0409_),
    .B(_0435_),
    .C(_0566_),
    .Y(\compressed_decoder_i.instr_o[1] ));
 sky130_fd_sc_hd__o21ai_0 _2161_ (.A1(\compressed_decoder_i.instr_i[2] ),
    .A2(_0455_),
    .B1(_0457_),
    .Y(_0567_));
 sky130_fd_sc_hd__nand2_1 _2162_ (.A(\compressed_decoder_i.instr_i[2] ),
    .B(_0444_),
    .Y(_0568_));
 sky130_fd_sc_hd__and2_0 _2163_ (.A(_0795_),
    .B(_0811_),
    .X(_0569_));
 sky130_fd_sc_hd__mux2_1 _2164_ (.A0(net170),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[20] ),
    .S(_0747_),
    .X(_0570_));
 sky130_fd_sc_hd__mux2i_4 _2165_ (.A0(_0570_),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[4] ),
    .S(_0836_),
    .Y(_0571_));
 sky130_fd_sc_hd__nor3_1 _2166_ (.A(_0434_),
    .B(_0519_),
    .C(_0571_),
    .Y(_0572_));
 sky130_fd_sc_hd__a31oi_1 _2167_ (.A1(\compressed_decoder_i.instr_i[15] ),
    .A2(_0519_),
    .A3(_0569_),
    .B1(_0572_),
    .Y(_0573_));
 sky130_fd_sc_hd__o21ai_0 _2168_ (.A1(_0411_),
    .A2(_0568_),
    .B1(_0573_),
    .Y(_0574_));
 sky130_fd_sc_hd__a21oi_1 _2169_ (.A1(_0447_),
    .A2(_0574_),
    .B1(_0540_),
    .Y(_0575_));
 sky130_fd_sc_hd__nand3_1 _2170_ (.A(\compressed_decoder_i.instr_i[2] ),
    .B(\compressed_decoder_i.instr_i[15] ),
    .C(_0488_),
    .Y(_0576_));
 sky130_fd_sc_hd__o21ai_0 _2171_ (.A1(_0533_),
    .A2(_0571_),
    .B1(_0576_),
    .Y(_0577_));
 sky130_fd_sc_hd__nor2_1 _2172_ (.A(\compressed_decoder_i.is_compressed_o ),
    .B(_0571_),
    .Y(_0578_));
 sky130_fd_sc_hd__a41oi_1 _2173_ (.A1(_0808_),
    .A2(_0414_),
    .A3(_0421_),
    .A4(_0459_),
    .B1(_0569_),
    .Y(_0579_));
 sky130_fd_sc_hd__a21oi_1 _2174_ (.A1(\compressed_decoder_i.instr_i[2] ),
    .A2(_0833_),
    .B1(_0791_),
    .Y(_0580_));
 sky130_fd_sc_hd__a221oi_1 _2175_ (.A1(\compressed_decoder_i.instr_i[13] ),
    .A2(_0571_),
    .B1(_0579_),
    .B2(_0580_),
    .C1(_0514_),
    .Y(_0581_));
 sky130_fd_sc_hd__a211oi_1 _2176_ (.A1(_0531_),
    .A2(_0577_),
    .B1(_0578_),
    .C1(_0581_),
    .Y(_0582_));
 sky130_fd_sc_hd__o21ai_1 _2177_ (.A1(_0567_),
    .A2(_0575_),
    .B1(_0582_),
    .Y(\compressed_decoder_i.instr_o[20] ));
 sky130_fd_sc_hd__mux2i_1 _2178_ (.A0(net171),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[21] ),
    .S(_0877_),
    .Y(_0583_));
 sky130_fd_sc_hd__nand2_1 _2179_ (.A(_0759_),
    .B(_0583_),
    .Y(_0584_));
 sky130_fd_sc_hd__o21ai_4 _2180_ (.A1(_0759_),
    .A2(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[5] ),
    .B1(_0584_),
    .Y(_0585_));
 sky130_fd_sc_hd__o22ai_1 _2181_ (.A1(_0475_),
    .A2(_0503_),
    .B1(_0519_),
    .B2(_0585_),
    .Y(_0586_));
 sky130_fd_sc_hd__nor2_2 _2182_ (.A(_0412_),
    .B(_0476_),
    .Y(_0587_));
 sky130_fd_sc_hd__a21oi_1 _2183_ (.A1(_0518_),
    .A2(_0586_),
    .B1(_0587_),
    .Y(_0588_));
 sky130_fd_sc_hd__and2_2 _2184_ (.A(\compressed_decoder_i.instr_o[0] ),
    .B(\compressed_decoder_i.is_compressed_o ),
    .X(_0589_));
 sky130_fd_sc_hd__o21ai_0 _2185_ (.A1(_0408_),
    .A2(_0798_),
    .B1(_0499_),
    .Y(_0590_));
 sky130_fd_sc_hd__a22oi_1 _2186_ (.A1(_0444_),
    .A2(_0456_),
    .B1(_0590_),
    .B2(_0468_),
    .Y(_0591_));
 sky130_fd_sc_hd__nor2_1 _2187_ (.A(\compressed_decoder_i.instr_i[13] ),
    .B(_0591_),
    .Y(_0592_));
 sky130_fd_sc_hd__a21oi_1 _2188_ (.A1(_0441_),
    .A2(_0501_),
    .B1(_0442_),
    .Y(_0593_));
 sky130_fd_sc_hd__o21ai_1 _2189_ (.A1(_0592_),
    .A2(_0593_),
    .B1(\compressed_decoder_i.instr_i[3] ),
    .Y(_0594_));
 sky130_fd_sc_hd__o221ai_4 _2190_ (.A1(_0458_),
    .A2(_0588_),
    .B1(_0589_),
    .B2(_0585_),
    .C1(_0594_),
    .Y(\compressed_decoder_i.instr_o[21] ));
 sky130_fd_sc_hd__clkinvlp_4 _2191_ (.A(\compressed_decoder_i.instr_i[4] ),
    .Y(_0595_));
 sky130_fd_sc_hd__mux2i_1 _2192_ (.A0(net172),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[22] ),
    .S(_0877_),
    .Y(_0596_));
 sky130_fd_sc_hd__nand2_1 _2193_ (.A(_0759_),
    .B(_0596_),
    .Y(_0597_));
 sky130_fd_sc_hd__o21ai_4 _2194_ (.A1(_0751_),
    .A2(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[6] ),
    .B1(_0597_),
    .Y(_0598_));
 sky130_fd_sc_hd__o22ai_1 _2195_ (.A1(_0595_),
    .A2(_0503_),
    .B1(_0519_),
    .B2(_0598_),
    .Y(_0599_));
 sky130_fd_sc_hd__o21ai_0 _2196_ (.A1(\compressed_decoder_i.instr_i[15] ),
    .A2(_0532_),
    .B1(_0501_),
    .Y(_0600_));
 sky130_fd_sc_hd__a221oi_2 _2197_ (.A1(_0518_),
    .A2(_0599_),
    .B1(_0600_),
    .B2(\compressed_decoder_i.instr_i[4] ),
    .C1(_0587_),
    .Y(_0601_));
 sky130_fd_sc_hd__nand2_2 _2198_ (.A(_0411_),
    .B(_0416_),
    .Y(_0602_));
 sky130_fd_sc_hd__nand2_1 _2199_ (.A(\compressed_decoder_i.instr_i[4] ),
    .B(_0457_),
    .Y(_0603_));
 sky130_fd_sc_hd__o22ai_1 _2200_ (.A1(\compressed_decoder_i.instr_i[6] ),
    .A2(\compressed_decoder_i.instr_i[15] ),
    .B1(_0499_),
    .B2(\compressed_decoder_i.instr_i[4] ),
    .Y(_0604_));
 sky130_fd_sc_hd__a22oi_1 _2201_ (.A1(_0595_),
    .A2(_0528_),
    .B1(_0604_),
    .B2(_0409_),
    .Y(_0605_));
 sky130_fd_sc_hd__a21oi_1 _2202_ (.A1(_0459_),
    .A2(_0598_),
    .B1(_0410_),
    .Y(_0606_));
 sky130_fd_sc_hd__nand2_1 _2203_ (.A(_0469_),
    .B(_0598_),
    .Y(_0607_));
 sky130_fd_sc_hd__o221ai_2 _2204_ (.A1(\compressed_decoder_i.instr_i[13] ),
    .A2(_0605_),
    .B1(_0606_),
    .B2(\compressed_decoder_i.instr_i[1] ),
    .C1(_0607_),
    .Y(_0608_));
 sky130_fd_sc_hd__o221ai_4 _2205_ (.A1(_0458_),
    .A2(_0601_),
    .B1(_0602_),
    .B2(_0603_),
    .C1(_0608_),
    .Y(\compressed_decoder_i.instr_o[22] ));
 sky130_fd_sc_hd__nor2b_1 _2206_ (.A(_0877_),
    .B_N(net173),
    .Y(_0609_));
 sky130_fd_sc_hd__a211oi_2 _2207_ (.A1(_0877_),
    .A2(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[23] ),
    .B1(_0609_),
    .C1(_0887_),
    .Y(_0610_));
 sky130_fd_sc_hd__a21oi_4 _2208_ (.A1(_0887_),
    .A2(_0824_),
    .B1(_0610_),
    .Y(_0611_));
 sky130_fd_sc_hd__nor2_1 _2209_ (.A(_0798_),
    .B(\compressed_decoder_i.instr_i[5] ),
    .Y(_0612_));
 sky130_fd_sc_hd__a21oi_1 _2210_ (.A1(\compressed_decoder_i.instr_i[14] ),
    .A2(_0548_),
    .B1(_0612_),
    .Y(_0613_));
 sky130_fd_sc_hd__o22ai_1 _2211_ (.A1(_0533_),
    .A2(_0611_),
    .B1(_0613_),
    .B2(_0431_),
    .Y(_0614_));
 sky130_fd_sc_hd__nor2_1 _2212_ (.A(_0512_),
    .B(_0460_),
    .Y(_0615_));
 sky130_fd_sc_hd__o21ai_0 _2213_ (.A1(_0412_),
    .A2(_0611_),
    .B1(_0615_),
    .Y(_0616_));
 sky130_fd_sc_hd__a22o_1 _2214_ (.A1(_0418_),
    .A2(_0488_),
    .B1(_0426_),
    .B2(_0460_),
    .X(_0617_));
 sky130_fd_sc_hd__nand2_1 _2215_ (.A(\compressed_decoder_i.instr_i[5] ),
    .B(_0617_),
    .Y(_0618_));
 sky130_fd_sc_hd__o211ai_1 _2216_ (.A1(_0412_),
    .A2(_0476_),
    .B1(_0616_),
    .C1(_0618_),
    .Y(_0619_));
 sky130_fd_sc_hd__a31oi_1 _2217_ (.A1(_0411_),
    .A2(\compressed_decoder_i.instr_i[5] ),
    .A3(_0416_),
    .B1(_0468_),
    .Y(_0620_));
 sky130_fd_sc_hd__nor2_1 _2218_ (.A(_0758_),
    .B(_0791_),
    .Y(_0621_));
 sky130_fd_sc_hd__nor2_1 _2219_ (.A(_0408_),
    .B(_0621_),
    .Y(_0622_));
 sky130_fd_sc_hd__a22oi_1 _2220_ (.A1(\compressed_decoder_i.instr_i[5] ),
    .A2(_0621_),
    .B1(_0622_),
    .B2(_0611_),
    .Y(_0623_));
 sky130_fd_sc_hd__o21ai_0 _2221_ (.A1(_0754_),
    .A2(_0620_),
    .B1(_0623_),
    .Y(_0624_));
 sky130_fd_sc_hd__a21oi_1 _2222_ (.A1(_0474_),
    .A2(_0619_),
    .B1(_0624_),
    .Y(_0625_));
 sky130_fd_sc_hd__a21oi_1 _2223_ (.A1(_0531_),
    .A2(_0614_),
    .B1(_0625_),
    .Y(\compressed_decoder_i.instr_o[23] ));
 sky130_fd_sc_hd__o21bai_1 _2224_ (.A1(_0464_),
    .A2(_0463_),
    .B1_N(_0617_),
    .Y(_0626_));
 sky130_fd_sc_hd__nor2_1 _2225_ (.A(_0751_),
    .B(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[8] ),
    .Y(_0627_));
 sky130_fd_sc_hd__nor2_1 _2226_ (.A(_0836_),
    .B(_0814_),
    .Y(_0628_));
 sky130_fd_sc_hd__nor2_2 _2227_ (.A(_0627_),
    .B(_0628_),
    .Y(_0629_));
 sky130_fd_sc_hd__a21oi_1 _2228_ (.A1(_0544_),
    .A2(_0629_),
    .B1(_0416_),
    .Y(_0630_));
 sky130_fd_sc_hd__a211oi_1 _2229_ (.A1(_0791_),
    .A2(_0424_),
    .B1(_0630_),
    .C1(_0798_),
    .Y(_0631_));
 sky130_fd_sc_hd__a311oi_1 _2230_ (.A1(\compressed_decoder_i.instr_i[6] ),
    .A2(_0457_),
    .A3(_0626_),
    .B1(_0631_),
    .C1(_0587_),
    .Y(_0632_));
 sky130_fd_sc_hd__o21ai_0 _2231_ (.A1(\compressed_decoder_i.instr_i[6] ),
    .A2(_0455_),
    .B1(_0457_),
    .Y(_0633_));
 sky130_fd_sc_hd__a221oi_1 _2232_ (.A1(\compressed_decoder_i.instr_i[11] ),
    .A2(_0452_),
    .B1(_0435_),
    .B2(_0629_),
    .C1(_0754_),
    .Y(_0634_));
 sky130_fd_sc_hd__a21oi_1 _2233_ (.A1(_0447_),
    .A2(\compressed_decoder_i.instr_i[6] ),
    .B1(_0409_),
    .Y(_0635_));
 sky130_fd_sc_hd__nor3_1 _2234_ (.A(_0410_),
    .B(_0634_),
    .C(_0635_),
    .Y(_0636_));
 sky130_fd_sc_hd__a21oi_1 _2235_ (.A1(_0622_),
    .A2(_0629_),
    .B1(_0636_),
    .Y(_0637_));
 sky130_fd_sc_hd__o21ai_0 _2236_ (.A1(_0632_),
    .A2(_0633_),
    .B1(_0637_),
    .Y(\compressed_decoder_i.instr_o[24] ));
 sky130_fd_sc_hd__o21ai_4 _2237_ (.A1(_0808_),
    .A2(_0455_),
    .B1(_0457_),
    .Y(_0638_));
 sky130_fd_sc_hd__nand3_1 _2238_ (.A(\compressed_decoder_i.instr_i[8] ),
    .B(_0420_),
    .C(_0429_),
    .Y(_0639_));
 sky130_fd_sc_hd__nor2_4 _2239_ (.A(_0485_),
    .B(_0538_),
    .Y(_0640_));
 sky130_fd_sc_hd__a21boi_0 _2240_ (.A1(_0639_),
    .A2(_0640_),
    .B1_N(\compressed_decoder_i.instr_i[2] ),
    .Y(_0641_));
 sky130_fd_sc_hd__nor2_1 _2241_ (.A(_0887_),
    .B(_0817_),
    .Y(_0642_));
 sky130_fd_sc_hd__a21oi_2 _2242_ (.A1(_0887_),
    .A2(_0825_),
    .B1(_0642_),
    .Y(_0643_));
 sky130_fd_sc_hd__nand3_2 _2243_ (.A(\compressed_decoder_i.instr_i[11] ),
    .B(_0808_),
    .C(_0426_),
    .Y(_0644_));
 sky130_fd_sc_hd__o21ba_1 _2244_ (.A1(_0548_),
    .A2(_0643_),
    .B1_N(_0644_),
    .X(_0645_));
 sky130_fd_sc_hd__a21oi_1 _2245_ (.A1(_0797_),
    .A2(_0463_),
    .B1(_0446_),
    .Y(_0646_));
 sky130_fd_sc_hd__a211oi_2 _2246_ (.A1(_0798_),
    .A2(_0806_),
    .B1(_0833_),
    .C1(_0646_),
    .Y(_0647_));
 sky130_fd_sc_hd__nor3_1 _2247_ (.A(_0641_),
    .B(_0645_),
    .C(_0647_),
    .Y(_0648_));
 sky130_fd_sc_hd__o21ai_0 _2248_ (.A1(_0754_),
    .A2(_0431_),
    .B1(_0532_),
    .Y(_0649_));
 sky130_fd_sc_hd__nand2_1 _2249_ (.A(\compressed_decoder_i.instr_o[0] ),
    .B(\compressed_decoder_i.is_compressed_o ),
    .Y(_0650_));
 sky130_fd_sc_hd__a32oi_1 _2250_ (.A1(_0468_),
    .A2(\compressed_decoder_i.instr_i[12] ),
    .A3(_0649_),
    .B1(_0643_),
    .B2(_0650_),
    .Y(_0651_));
 sky130_fd_sc_hd__o21ai_1 _2251_ (.A1(_0638_),
    .A2(_0648_),
    .B1(_0651_),
    .Y(\compressed_decoder_i.instr_o[25] ));
 sky130_fd_sc_hd__mux2i_1 _2252_ (.A0(net176),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[26] ),
    .S(_0877_),
    .Y(_0652_));
 sky130_fd_sc_hd__nand2_1 _2253_ (.A(_0759_),
    .B(_0652_),
    .Y(_0653_));
 sky130_fd_sc_hd__o21ai_2 _2254_ (.A1(_0751_),
    .A2(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[10] ),
    .B1(_0653_),
    .Y(_0654_));
 sky130_fd_sc_hd__a21oi_1 _2255_ (.A1(\compressed_decoder_i.instr_i[10] ),
    .A2(_0654_),
    .B1(_0644_),
    .Y(_0655_));
 sky130_fd_sc_hd__a21boi_0 _2256_ (.A1(_0499_),
    .A2(_0639_),
    .B1_N(\compressed_decoder_i.instr_i[5] ),
    .Y(_0656_));
 sky130_fd_sc_hd__a2111oi_0 _2257_ (.A1(\compressed_decoder_i.instr_i[7] ),
    .A2(_0485_),
    .B1(_0647_),
    .C1(_0655_),
    .D1(_0656_),
    .Y(_0657_));
 sky130_fd_sc_hd__nand2_1 _2258_ (.A(_0435_),
    .B(_0654_),
    .Y(_0658_));
 sky130_fd_sc_hd__o221ai_1 _2259_ (.A1(\compressed_decoder_i.instr_i[5] ),
    .A2(_0532_),
    .B1(_0455_),
    .B2(\compressed_decoder_i.instr_i[7] ),
    .C1(_0531_),
    .Y(_0659_));
 sky130_fd_sc_hd__o21ai_0 _2260_ (.A1(_0551_),
    .A2(_0654_),
    .B1(_0659_),
    .Y(_0660_));
 sky130_fd_sc_hd__nand2_1 _2261_ (.A(\compressed_decoder_i.instr_i[7] ),
    .B(\compressed_decoder_i.instr_i[15] ),
    .Y(_0661_));
 sky130_fd_sc_hd__a211oi_2 _2262_ (.A1(_0568_),
    .A2(_0661_),
    .B1(_0532_),
    .C1(_0514_),
    .Y(_0662_));
 sky130_fd_sc_hd__a21oi_1 _2263_ (.A1(_0658_),
    .A2(_0660_),
    .B1(_0662_),
    .Y(_0663_));
 sky130_fd_sc_hd__o21ai_1 _2264_ (.A1(_0638_),
    .A2(_0657_),
    .B1(_0663_),
    .Y(\compressed_decoder_i.instr_o[26] ));
 sky130_fd_sc_hd__nor2_1 _2265_ (.A(_0477_),
    .B(_0640_),
    .Y(_0664_));
 sky130_fd_sc_hd__mux2i_1 _2266_ (.A0(net177),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[27] ),
    .S(_0877_),
    .Y(_0665_));
 sky130_fd_sc_hd__nand2_1 _2267_ (.A(_0759_),
    .B(_0665_),
    .Y(_0666_));
 sky130_fd_sc_hd__o21ai_2 _2268_ (.A1(_0759_),
    .A2(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[11] ),
    .B1(_0666_),
    .Y(_0667_));
 sky130_fd_sc_hd__a21oi_1 _2269_ (.A1(\compressed_decoder_i.instr_i[10] ),
    .A2(_0667_),
    .B1(_0644_),
    .Y(_0668_));
 sky130_fd_sc_hd__a2111oi_0 _2270_ (.A1(\compressed_decoder_i.instr_i[3] ),
    .A2(_0525_),
    .B1(_0647_),
    .C1(_0664_),
    .D1(_0668_),
    .Y(_0669_));
 sky130_fd_sc_hd__nand2_1 _2271_ (.A(_0816_),
    .B(_0432_),
    .Y(_0670_));
 sky130_fd_sc_hd__nand2_1 _2272_ (.A(_0431_),
    .B(_0667_),
    .Y(_0671_));
 sky130_fd_sc_hd__nor2_1 _2273_ (.A(_0816_),
    .B(_0418_),
    .Y(_0672_));
 sky130_fd_sc_hd__a21oi_1 _2274_ (.A1(\compressed_decoder_i.instr_i[3] ),
    .A2(_0444_),
    .B1(_0672_),
    .Y(_0673_));
 sky130_fd_sc_hd__o32ai_1 _2275_ (.A1(_0532_),
    .A2(_0514_),
    .A3(_0673_),
    .B1(_0667_),
    .B2(_0551_),
    .Y(_0674_));
 sky130_fd_sc_hd__a31oi_1 _2276_ (.A1(_0670_),
    .A2(_0554_),
    .A3(_0671_),
    .B1(_0674_),
    .Y(_0675_));
 sky130_fd_sc_hd__o21ai_0 _2277_ (.A1(_0638_),
    .A2(_0669_),
    .B1(_0675_),
    .Y(\compressed_decoder_i.instr_o[27] ));
 sky130_fd_sc_hd__nand2_1 _2278_ (.A(_0887_),
    .B(_0827_),
    .Y(_0676_));
 sky130_fd_sc_hd__o21ai_2 _2279_ (.A1(_0836_),
    .A2(_0804_),
    .B1(_0676_),
    .Y(_0677_));
 sky130_fd_sc_hd__o22ai_1 _2280_ (.A1(_0820_),
    .A2(_0441_),
    .B1(_0499_),
    .B2(_0806_),
    .Y(_0678_));
 sky130_fd_sc_hd__a21oi_1 _2281_ (.A1(\compressed_decoder_i.instr_i[10] ),
    .A2(_0677_),
    .B1(_0644_),
    .Y(_0679_));
 sky130_fd_sc_hd__a2111oi_0 _2282_ (.A1(\compressed_decoder_i.instr_i[4] ),
    .A2(_0525_),
    .B1(_0647_),
    .C1(_0678_),
    .D1(_0679_),
    .Y(_0680_));
 sky130_fd_sc_hd__nand2_1 _2283_ (.A(_0431_),
    .B(_0677_),
    .Y(_0681_));
 sky130_fd_sc_hd__nand3_1 _2284_ (.A(_0542_),
    .B(_0554_),
    .C(_0681_),
    .Y(_0682_));
 sky130_fd_sc_hd__o221ai_1 _2285_ (.A1(_0551_),
    .A2(_0677_),
    .B1(_0680_),
    .B2(_0638_),
    .C1(_0682_),
    .Y(\compressed_decoder_i.instr_o[28] ));
 sky130_fd_sc_hd__nand2_1 _2286_ (.A(_0887_),
    .B(_0828_),
    .Y(_0683_));
 sky130_fd_sc_hd__o21ai_2 _2287_ (.A1(_0887_),
    .A2(_0786_),
    .B1(_0683_),
    .Y(_0684_));
 sky130_fd_sc_hd__a21oi_1 _2288_ (.A1(_0791_),
    .A2(_0548_),
    .B1(_0602_),
    .Y(_0685_));
 sky130_fd_sc_hd__a21oi_1 _2289_ (.A1(\compressed_decoder_i.instr_i[10] ),
    .A2(_0684_),
    .B1(_0644_),
    .Y(_0686_));
 sky130_fd_sc_hd__a211oi_1 _2290_ (.A1(\compressed_decoder_i.instr_i[14] ),
    .A2(\compressed_decoder_i.instr_i[12] ),
    .B1(_0685_),
    .C1(_0686_),
    .Y(_0687_));
 sky130_fd_sc_hd__nand2_1 _2291_ (.A(_0431_),
    .B(_0684_),
    .Y(_0688_));
 sky130_fd_sc_hd__nand3_1 _2292_ (.A(_0549_),
    .B(_0554_),
    .C(_0688_),
    .Y(_0689_));
 sky130_fd_sc_hd__o221ai_1 _2293_ (.A1(_0551_),
    .A2(_0684_),
    .B1(_0687_),
    .B2(_0638_),
    .C1(_0689_),
    .Y(\compressed_decoder_i.instr_o[29] ));
 sky130_fd_sc_hd__nand2_1 _2294_ (.A(_0808_),
    .B(_0421_),
    .Y(_0690_));
 sky130_fd_sc_hd__nand3_1 _2295_ (.A(_0447_),
    .B(_0415_),
    .C(_0690_),
    .Y(_0691_));
 sky130_fd_sc_hd__a2bb2oi_1 _2296_ (.A1_N(_0434_),
    .A2_N(_0691_),
    .B1(\compressed_decoder_i.instr_i[13] ),
    .B2(\compressed_decoder_i.instr_i[2] ),
    .Y(_0692_));
 sky130_fd_sc_hd__a21oi_1 _2297_ (.A1(_0441_),
    .A2(_0476_),
    .B1(_0458_),
    .Y(_0693_));
 sky130_fd_sc_hd__a21oi_1 _2298_ (.A1(\compressed_decoder_i.instr_i[2] ),
    .A2(_0564_),
    .B1(_0693_),
    .Y(_0694_));
 sky130_fd_sc_hd__o21ai_0 _2299_ (.A1(_0514_),
    .A2(_0692_),
    .B1(_0694_),
    .Y(\compressed_decoder_i.instr_o[2] ));
 sky130_fd_sc_hd__mux2i_4 _2300_ (.A0(_0792_),
    .A1(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[14] ),
    .S(_0836_),
    .Y(_0695_));
 sky130_fd_sc_hd__nand2_1 _2301_ (.A(_0801_),
    .B(_0695_),
    .Y(_0696_));
 sky130_fd_sc_hd__a31oi_1 _2302_ (.A1(\compressed_decoder_i.instr_i[11] ),
    .A2(_0808_),
    .A3(_0696_),
    .B1(_0416_),
    .Y(_0697_));
 sky130_fd_sc_hd__o21ai_0 _2303_ (.A1(_0424_),
    .A2(_0433_),
    .B1(\compressed_decoder_i.instr_i[10] ),
    .Y(_0698_));
 sky130_fd_sc_hd__a221oi_1 _2304_ (.A1(_0791_),
    .A2(_0816_),
    .B1(_0697_),
    .B2(_0698_),
    .C1(\compressed_decoder_i.instr_i[14] ),
    .Y(_0699_));
 sky130_fd_sc_hd__a21oi_1 _2305_ (.A1(\compressed_decoder_i.instr_i[14] ),
    .A2(\compressed_decoder_i.instr_i[12] ),
    .B1(_0699_),
    .Y(_0700_));
 sky130_fd_sc_hd__o22ai_1 _2306_ (.A1(_0589_),
    .A2(_0695_),
    .B1(_0700_),
    .B2(_0638_),
    .Y(\compressed_decoder_i.instr_o[30] ));
 sky130_fd_sc_hd__mux2i_4 _2307_ (.A0(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[15] ),
    .A1(_0829_),
    .S(_0759_),
    .Y(_0701_));
 sky130_fd_sc_hd__nand2_1 _2308_ (.A(\compressed_decoder_i.instr_i[10] ),
    .B(_0701_),
    .Y(_0702_));
 sky130_fd_sc_hd__a21oi_1 _2309_ (.A1(\compressed_decoder_i.instr_i[11] ),
    .A2(_0702_),
    .B1(_0512_),
    .Y(_0703_));
 sky130_fd_sc_hd__o32ai_2 _2310_ (.A1(_0412_),
    .A2(_0442_),
    .A3(_0703_),
    .B1(_0701_),
    .B2(_0589_),
    .Y(\compressed_decoder_i.instr_o[31] ));
 sky130_fd_sc_hd__a31oi_1 _2311_ (.A1(_0459_),
    .A2(_0474_),
    .A3(_0544_),
    .B1(_0650_),
    .Y(_0704_));
 sky130_fd_sc_hd__o22ai_1 _2312_ (.A1(_0441_),
    .A2(_0442_),
    .B1(_0704_),
    .B2(_0475_),
    .Y(\compressed_decoder_i.instr_o[3] ));
 sky130_fd_sc_hd__o21ai_0 _2313_ (.A1(_0754_),
    .A2(_0444_),
    .B1(_0446_),
    .Y(_0705_));
 sky130_fd_sc_hd__a21oi_1 _2314_ (.A1(_0595_),
    .A2(_0705_),
    .B1(_0488_),
    .Y(_0706_));
 sky130_fd_sc_hd__o31ai_1 _2315_ (.A1(_0409_),
    .A2(_0444_),
    .A3(_0691_),
    .B1(_0706_),
    .Y(_0707_));
 sky130_fd_sc_hd__a21oi_1 _2316_ (.A1(\compressed_decoder_i.instr_i[15] ),
    .A2(_0544_),
    .B1(_0754_),
    .Y(_0708_));
 sky130_fd_sc_hd__o221ai_1 _2317_ (.A1(\compressed_decoder_i.instr_i[1] ),
    .A2(_0640_),
    .B1(_0708_),
    .B2(\compressed_decoder_i.instr_i[4] ),
    .C1(\compressed_decoder_i.instr_i[0] ),
    .Y(_0709_));
 sky130_fd_sc_hd__o21ai_1 _2318_ (.A1(\compressed_decoder_i.instr_i[0] ),
    .A2(_0707_),
    .B1(_0709_),
    .Y(\compressed_decoder_i.instr_o[4] ));
 sky130_fd_sc_hd__o21ai_0 _2319_ (.A1(\compressed_decoder_i.instr_i[5] ),
    .A2(_0806_),
    .B1(_0615_),
    .Y(_0710_));
 sky130_fd_sc_hd__and3_1 _2320_ (.A(_0476_),
    .B(_0640_),
    .C(_0710_),
    .X(_0711_));
 sky130_fd_sc_hd__o21ai_0 _2321_ (.A1(_0410_),
    .A2(_0612_),
    .B1(_0409_),
    .Y(_0712_));
 sky130_fd_sc_hd__o221ai_1 _2322_ (.A1(_0410_),
    .A2(_0431_),
    .B1(_0621_),
    .B2(\compressed_decoder_i.instr_i[5] ),
    .C1(_0712_),
    .Y(_0713_));
 sky130_fd_sc_hd__o21ai_0 _2323_ (.A1(_0458_),
    .A2(_0711_),
    .B1(_0713_),
    .Y(\compressed_decoder_i.instr_o[5] ));
 sky130_fd_sc_hd__a21oi_1 _2324_ (.A1(\compressed_decoder_i.instr_i[13] ),
    .A2(_0528_),
    .B1(_0564_),
    .Y(_0714_));
 sky130_fd_sc_hd__nand4_1 _2325_ (.A(\compressed_decoder_i.instr_i[1] ),
    .B(_0468_),
    .C(_0415_),
    .D(_0426_),
    .Y(_0715_));
 sky130_fd_sc_hd__o221ai_2 _2326_ (.A1(_0442_),
    .A2(_0640_),
    .B1(_0714_),
    .B2(_0477_),
    .C1(_0715_),
    .Y(\compressed_decoder_i.instr_o[6] ));
 sky130_fd_sc_hd__o21ai_0 _2327_ (.A1(_0412_),
    .A2(_0421_),
    .B1(_0415_),
    .Y(_0716_));
 sky130_fd_sc_hd__a211oi_1 _2328_ (.A1(_0411_),
    .A2(_0716_),
    .B1(_0514_),
    .C1(_0416_),
    .Y(_0717_));
 sky130_fd_sc_hd__nor4_1 _2329_ (.A(\compressed_decoder_i.instr_i[7] ),
    .B(_0444_),
    .C(_0415_),
    .D(_0514_),
    .Y(_0718_));
 sky130_fd_sc_hd__a21oi_1 _2330_ (.A1(_0757_),
    .A2(_0426_),
    .B1(_0408_),
    .Y(_0719_));
 sky130_fd_sc_hd__a21oi_1 _2331_ (.A1(_0410_),
    .A2(_0432_),
    .B1(_0719_),
    .Y(_0720_));
 sky130_fd_sc_hd__a21oi_1 _2332_ (.A1(\compressed_decoder_i.instr_i[2] ),
    .A2(_0452_),
    .B1(_0510_),
    .Y(_0721_));
 sky130_fd_sc_hd__o21ai_1 _2333_ (.A1(_0492_),
    .A2(_0533_),
    .B1(_0721_),
    .Y(_0722_));
 sky130_fd_sc_hd__a21oi_1 _2334_ (.A1(_0446_),
    .A2(\compressed_decoder_i.instr_i[7] ),
    .B1(_0444_),
    .Y(_0723_));
 sky130_fd_sc_hd__a221oi_1 _2335_ (.A1(\compressed_decoder_i.instr_i[7] ),
    .A2(_0418_),
    .B1(_0538_),
    .B2(_0808_),
    .C1(_0442_),
    .Y(_0724_));
 sky130_fd_sc_hd__o21ai_0 _2336_ (.A1(\compressed_decoder_i.instr_i[14] ),
    .A2(_0723_),
    .B1(_0724_),
    .Y(_0725_));
 sky130_fd_sc_hd__o211ai_2 _2337_ (.A1(\compressed_decoder_i.instr_i[7] ),
    .A2(_0720_),
    .B1(_0722_),
    .C1(_0725_),
    .Y(_0726_));
 sky130_fd_sc_hd__nor3_1 _2338_ (.A(_0717_),
    .B(_0718_),
    .C(_0726_),
    .Y(\compressed_decoder_i.instr_o[7] ));
 sky130_fd_sc_hd__a22oi_1 _2339_ (.A1(\compressed_decoder_i.instr_i[3] ),
    .A2(_0452_),
    .B1(_0435_),
    .B2(\compressed_decoder_i.instr_i[8] ),
    .Y(_0727_));
 sky130_fd_sc_hd__nor2_1 _2340_ (.A(\compressed_decoder_i.instr_i[14] ),
    .B(_0415_),
    .Y(_0728_));
 sky130_fd_sc_hd__nor3_1 _2341_ (.A(\compressed_decoder_i.instr_i[0] ),
    .B(_0416_),
    .C(_0728_),
    .Y(_0729_));
 sky130_fd_sc_hd__nand3_1 _2342_ (.A(_0408_),
    .B(\compressed_decoder_i.instr_i[3] ),
    .C(_0538_),
    .Y(_0730_));
 sky130_fd_sc_hd__o21ai_0 _2343_ (.A1(_0816_),
    .A2(_0538_),
    .B1(_0730_),
    .Y(_0731_));
 sky130_fd_sc_hd__a32oi_1 _2344_ (.A1(\compressed_decoder_i.instr_i[0] ),
    .A2(_0441_),
    .A3(_0731_),
    .B1(\compressed_decoder_i.instr_i[8] ),
    .B2(\compressed_decoder_i.instr_i[1] ),
    .Y(_0732_));
 sky130_fd_sc_hd__o22ai_1 _2345_ (.A1(_0510_),
    .A2(_0727_),
    .B1(_0729_),
    .B2(_0732_),
    .Y(\compressed_decoder_i.instr_o[8] ));
 sky130_fd_sc_hd__o21ai_0 _2346_ (.A1(\compressed_decoder_i.instr_i[9] ),
    .A2(_0418_),
    .B1(_0446_),
    .Y(_0733_));
 sky130_fd_sc_hd__nor2_1 _2347_ (.A(\compressed_decoder_i.instr_i[9] ),
    .B(_0833_),
    .Y(_0734_));
 sky130_fd_sc_hd__a21oi_1 _2348_ (.A1(_0595_),
    .A2(_0833_),
    .B1(_0734_),
    .Y(_0735_));
 sky130_fd_sc_hd__nor2_1 _2349_ (.A(_0411_),
    .B(_0735_),
    .Y(_0736_));
 sky130_fd_sc_hd__a21oi_1 _2350_ (.A1(_0411_),
    .A2(_0733_),
    .B1(_0736_),
    .Y(_0737_));
 sky130_fd_sc_hd__a31oi_1 _2351_ (.A1(_0468_),
    .A2(_0415_),
    .A3(_0426_),
    .B1(_0409_),
    .Y(_0738_));
 sky130_fd_sc_hd__a21oi_1 _2352_ (.A1(\compressed_decoder_i.instr_i[0] ),
    .A2(_0737_),
    .B1(_0738_),
    .Y(_0739_));
 sky130_fd_sc_hd__nand3_1 _2353_ (.A(_0798_),
    .B(_0477_),
    .C(_0833_),
    .Y(_0740_));
 sky130_fd_sc_hd__o21ai_0 _2354_ (.A1(\compressed_decoder_i.instr_i[4] ),
    .A2(\compressed_decoder_i.instr_i[15] ),
    .B1(_0740_),
    .Y(_0741_));
 sky130_fd_sc_hd__a221oi_1 _2355_ (.A1(_0820_),
    .A2(_0435_),
    .B1(_0741_),
    .B2(_0447_),
    .C1(_0510_),
    .Y(_0742_));
 sky130_fd_sc_hd__a21oi_1 _2356_ (.A1(_0474_),
    .A2(_0737_),
    .B1(_0742_),
    .Y(_0743_));
 sky130_fd_sc_hd__o21ai_1 _2357_ (.A1(_0820_),
    .A2(_0739_),
    .B1(_0743_),
    .Y(\compressed_decoder_i.instr_o[9] ));
 sky130_fd_sc_hd__inv_1 _2358_ (.A(net316),
    .Y(_0744_));
 sky130_fd_sc_hd__o22ai_1 _2359_ (.A1(_0744_),
    .A2(net191),
    .B1(_0785_),
    .B2(_0844_),
    .Y(instr_valid_id_d));
 sky130_fd_sc_hd__fa_1 _2360_ (.A(net369),
    .B(_1056_),
    .CIN(_1057_),
    .COUT(_1058_),
    .SUM(_1059_));
 sky130_fd_sc_hd__ha_1 _2361_ (.A(net358),
    .B(_1060_),
    .COUT(_1056_),
    .SUM(_1061_));
 sky130_fd_sc_hd__ha_1 _2362_ (.A(net369),
    .B(_1057_),
    .COUT(_1062_),
    .SUM(_1063_));
 sky130_fd_sc_hd__ha_1 _2363_ (.A(_1064_),
    .B(_1065_),
    .COUT(_1066_),
    .SUM(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[2] ));
 sky130_fd_sc_hd__ha_1 _2364_ (.A(_1067_),
    .B(_1066_),
    .COUT(_1068_),
    .SUM(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[3] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk_i (.A(clknet_2_0__leaf_clk_i),
    .X(clknet_leaf_0_clk_i));
 sky130_fd_sc_hd__buf_4 _2366_ (.A(net379),
    .X(dummy_instr_id_o));
 sky130_fd_sc_hd__buf_4 _2367_ (.A(net380),
    .X(instr_addr_o[0]));
 sky130_fd_sc_hd__buf_4 _2368_ (.A(net381),
    .X(instr_addr_o[1]));
 sky130_fd_sc_hd__buf_4 _2369_ (.A(net382),
    .X(instr_bp_taken_o));
 sky130_fd_sc_hd__clkbuf_1 _2370_ (.A(net235),
    .X(net283));
 sky130_fd_sc_hd__clkbuf_2 _2371_ (.A(net246),
    .X(net294));
 sky130_fd_sc_hd__clkbuf_1 _2372_ (.A(net257),
    .X(net305));
 sky130_fd_sc_hd__clkbuf_2 _2373_ (.A(net260),
    .X(net308));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2374_ (.A(net261),
    .X(net309));
 sky130_fd_sc_hd__clkbuf_1 _2375_ (.A(net262),
    .X(net310));
 sky130_fd_sc_hd__clkbuf_1 _2376_ (.A(net263),
    .X(net311));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2377_ (.A(net264),
    .X(net312));
 sky130_fd_sc_hd__clkbuf_1 _2378_ (.A(net265),
    .X(net313));
 sky130_fd_sc_hd__clkbuf_2 _2379_ (.A(net266),
    .X(net314));
 sky130_fd_sc_hd__clkbuf_1 _2380_ (.A(net236),
    .X(net284));
 sky130_fd_sc_hd__clkbuf_1 _2381_ (.A(net237),
    .X(net285));
 sky130_fd_sc_hd__clkbuf_2 _2382_ (.A(net238),
    .X(net286));
 sky130_fd_sc_hd__clkbuf_2 _2383_ (.A(net239),
    .X(net287));
 sky130_fd_sc_hd__buf_2 _2384_ (.A(net240),
    .X(net288));
 sky130_fd_sc_hd__clkbuf_1 _2385_ (.A(net241),
    .X(net289));
 sky130_fd_sc_hd__buf_2 _2386_ (.A(net242),
    .X(net290));
 sky130_fd_sc_hd__clkbuf_2 _2387_ (.A(net243),
    .X(net291));
 sky130_fd_sc_hd__clkbuf_1 _2388_ (.A(net244),
    .X(net292));
 sky130_fd_sc_hd__clkbuf_1 _2389_ (.A(net245),
    .X(net293));
 sky130_fd_sc_hd__clkbuf_2 _2390_ (.A(net247),
    .X(net295));
 sky130_fd_sc_hd__clkbuf_1 _2391_ (.A(net248),
    .X(net296));
 sky130_fd_sc_hd__clkbuf_1 _2392_ (.A(net249),
    .X(net297));
 sky130_fd_sc_hd__clkbuf_1 _2393_ (.A(net250),
    .X(net298));
 sky130_fd_sc_hd__clkbuf_1 _2394_ (.A(net251),
    .X(net299));
 sky130_fd_sc_hd__clkbuf_1 _2395_ (.A(net252),
    .X(net300));
 sky130_fd_sc_hd__clkbuf_1 _2396_ (.A(net253),
    .X(net301));
 sky130_fd_sc_hd__clkbuf_1 _2397_ (.A(net254),
    .X(net302));
 sky130_fd_sc_hd__clkbuf_1 _2398_ (.A(net255),
    .X(net303));
 sky130_fd_sc_hd__clkbuf_1 _2399_ (.A(net256),
    .X(net304));
 sky130_fd_sc_hd__clkbuf_1 _2400_ (.A(net258),
    .X(net306));
 sky130_fd_sc_hd__clkbuf_1 _2401_ (.A(net259),
    .X(net307));
 sky130_fd_sc_hd__buf_4 _2402_ (.A(net383),
    .X(pc_id_o[0]));
 sky130_fd_sc_hd__buf_4 _2403_ (.A(net384),
    .X(pc_if_o[0]));
 sky130_fd_sc_hd__buf_4 _2404_ (.A(net385),
    .X(pc_mismatch_alert_o));
 sky130_fd_sc_hd__dfrtp_4 \gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0]$_DFF_PN0_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[0] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[0] ),
    .RESET_B(net197),
    .CLK(clknet_leaf_30_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[1]$_DFF_PN0_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.branch_discard_s[1] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.branch_discard_q[1] ),
    .RESET_B(net197),
    .CLK(clknet_leaf_30_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \gen_prefetch_buffer.prefetch_buffer_i.discard_req_q$_DFF_PN0_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.discard_req_d ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.discard_req_q ),
    .RESET_B(net197),
    .CLK(clknet_leaf_34_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[10]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[10] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[10] ),
    .CLK(clknet_leaf_3_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[11]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[11] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[11] ),
    .CLK(clknet_leaf_2_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[12]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[12] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[12] ),
    .CLK(clknet_leaf_3_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[13]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[13] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[13] ),
    .CLK(clknet_leaf_3_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[14]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[14] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[14] ),
    .CLK(clknet_leaf_3_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[15]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[15] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[15] ),
    .CLK(clknet_leaf_2_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[16]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[16] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[16] ),
    .CLK(clknet_leaf_2_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[17]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[17] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[17] ),
    .CLK(clknet_leaf_33_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[18]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[18] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[18] ),
    .CLK(clknet_leaf_3_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[19]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[19] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[19] ),
    .CLK(clknet_leaf_32_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[20]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[20] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[20] ),
    .CLK(clknet_leaf_32_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[21]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[21] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[21] ),
    .CLK(clknet_leaf_3_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[22]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[22] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[22] ),
    .CLK(clknet_leaf_3_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[23]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[23] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[23] ),
    .CLK(clknet_leaf_4_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[24]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[24] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[24] ),
    .CLK(clknet_leaf_4_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[25]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[25] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[25] ),
    .CLK(clknet_leaf_4_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[26]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[26] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[26] ),
    .CLK(clknet_leaf_4_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[27]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[27] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[27] ),
    .CLK(clknet_leaf_4_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[28]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[28] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[28] ),
    .CLK(clknet_leaf_4_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[29]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[29] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[29] ),
    .CLK(clknet_leaf_4_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[2]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[2] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[2] ),
    .CLK(clknet_leaf_0_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[30]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[30] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[30] ),
    .CLK(clknet_leaf_3_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[31]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[31] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[31] ),
    .CLK(clknet_leaf_8_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[3]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[3] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[3] ),
    .CLK(clknet_leaf_1_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[4]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[4] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[4] ),
    .CLK(clknet_leaf_1_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[5]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[5] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[5] ),
    .CLK(clknet_leaf_1_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[6]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[6] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[6] ),
    .CLK(clknet_leaf_1_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[7]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[7] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[7] ),
    .CLK(clknet_leaf_1_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[8]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[8] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[8] ),
    .CLK(clknet_leaf_1_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[9]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_d[9] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fetch_addr_q[9] ),
    .CLK(clknet_leaf_2_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[0]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_d[0] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[0] ),
    .CLK(clknet_leaf_31_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_d[1] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[1] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[1] ),
    .CLK(clknet_leaf_31_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[2]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_d[2] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[2] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.err_q[2] ),
    .CLK(clknet_leaf_31_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[0]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[1] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_en ),
    .Q(net358),
    .CLK(clknet_leaf_1_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[10]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[11] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_en ),
    .Q(net349),
    .CLK(clknet_leaf_11_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[11]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[12] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_en ),
    .Q(net350),
    .CLK(clknet_leaf_11_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[12]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[13] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_en ),
    .Q(net351),
    .CLK(clknet_leaf_9_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[13]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[14] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_en ),
    .Q(net352),
    .CLK(clknet_leaf_8_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[14]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[15] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_en ),
    .Q(net353),
    .CLK(clknet_leaf_8_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[15]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[16] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_en ),
    .Q(net354),
    .CLK(clknet_leaf_9_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[16]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[17] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_en ),
    .Q(net355),
    .CLK(clknet_leaf_7_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[17]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[18] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_en ),
    .Q(net356),
    .CLK(clknet_leaf_7_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[18]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[19] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_en ),
    .Q(net357),
    .CLK(clknet_leaf_7_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[19]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[20] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_en ),
    .Q(net359),
    .CLK(clknet_leaf_7_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[1]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[2] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_en ),
    .Q(net369),
    .CLK(clknet_leaf_1_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[20]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[21] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_en ),
    .Q(net360),
    .CLK(clknet_leaf_7_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[21]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[22] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_en ),
    .Q(net361),
    .CLK(clknet_leaf_11_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[22]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[23] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_en ),
    .Q(net362),
    .CLK(clknet_leaf_6_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[23]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[24] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_en ),
    .Q(net363),
    .CLK(clknet_leaf_12_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[24]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[25] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_en ),
    .Q(net364),
    .CLK(clknet_leaf_6_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[25]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[26] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_en ),
    .Q(net365),
    .CLK(clknet_leaf_11_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[26]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[27] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_en ),
    .Q(net366),
    .CLK(clknet_leaf_11_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[27]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[28] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_en ),
    .Q(net367),
    .CLK(clknet_leaf_6_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[28]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[29] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_en ),
    .Q(net368),
    .CLK(clknet_leaf_6_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[29]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[30] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_en ),
    .Q(net370),
    .CLK(clknet_leaf_6_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[2]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[3] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_en ),
    .Q(net372),
    .CLK(clknet_leaf_8_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[30]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[31] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_en ),
    .Q(net371),
    .CLK(clknet_leaf_7_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[3]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[4] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_en ),
    .Q(net373),
    .CLK(clknet_leaf_9_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[4]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[5] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_en ),
    .Q(net374),
    .CLK(clknet_leaf_8_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[5]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[6] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_en ),
    .Q(net375),
    .CLK(clknet_leaf_8_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[6]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[7] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_en ),
    .Q(net376),
    .CLK(clknet_leaf_9_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[7]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[8] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_en ),
    .Q(net377),
    .CLK(clknet_leaf_8_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[8]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[9] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_en ),
    .Q(net378),
    .CLK(clknet_leaf_9_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_q[9]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_d[10] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.instr_addr_en ),
    .Q(net348),
    .CLK(clknet_leaf_11_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[0]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[0] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[0] ),
    .CLK(clknet_leaf_29_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[10]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[10] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[10] ),
    .CLK(clknet_leaf_24_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[11]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[11] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[11] ),
    .CLK(clknet_leaf_24_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[12]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[12] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[12] ),
    .CLK(clknet_leaf_20_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[13]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[13] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[13] ),
    .CLK(clknet_leaf_21_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[14]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[14] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[14] ),
    .CLK(clknet_leaf_18_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[15]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[15] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[15] ),
    .CLK(clknet_leaf_20_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[16]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[16] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[16] ),
    .CLK(clknet_leaf_27_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[17]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[17] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[17] ),
    .CLK(clknet_leaf_31_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[18]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[18] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[18] ),
    .CLK(clknet_leaf_26_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[19]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[19] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[19] ),
    .CLK(clknet_leaf_26_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[1]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[1] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[1] ),
    .CLK(clknet_leaf_29_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[20]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[20] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[20] ),
    .CLK(clknet_leaf_27_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[21]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[21] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[21] ),
    .CLK(clknet_leaf_26_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[22]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[22] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[22] ),
    .CLK(clknet_leaf_28_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[23]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[23] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[23] ),
    .CLK(clknet_leaf_24_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[24]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[24] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[24] ),
    .CLK(clknet_leaf_25_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[25]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[25] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[25] ),
    .CLK(clknet_leaf_23_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[26]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[26] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[26] ),
    .CLK(clknet_leaf_25_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[27]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[27] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[27] ),
    .CLK(clknet_leaf_24_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[28]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[28] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[28] ),
    .CLK(clknet_leaf_22_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[29]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[29] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[29] ),
    .CLK(clknet_leaf_22_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[2]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[2] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[2] ),
    .CLK(clknet_leaf_28_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[30]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[30] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[30] ),
    .CLK(clknet_leaf_23_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[31]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[31] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[31] ),
    .CLK(clknet_leaf_22_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[32]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[32] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[1] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[32] ),
    .CLK(clknet_leaf_30_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[33]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[33] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[1] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[33] ),
    .CLK(clknet_leaf_29_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[34]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[34] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[1] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[34] ),
    .CLK(clknet_leaf_28_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[35]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[35] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[1] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[35] ),
    .CLK(clknet_leaf_27_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[36]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[36] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[1] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[36] ),
    .CLK(clknet_leaf_29_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[37]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[37] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[1] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[37] ),
    .CLK(clknet_leaf_25_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[38]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[38] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[1] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[38] ),
    .CLK(clknet_leaf_28_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[39]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[39] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[1] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[39] ),
    .CLK(clknet_leaf_22_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[3]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[3] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[3] ),
    .CLK(clknet_leaf_27_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[40]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[40] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[1] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[40] ),
    .CLK(clknet_leaf_28_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[41]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[41] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[1] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[41] ),
    .CLK(clknet_leaf_20_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[42]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[42] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[1] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[42] ),
    .CLK(clknet_leaf_24_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[43]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[43] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[1] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[43] ),
    .CLK(clknet_leaf_21_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[44]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[44] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[1] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[44] ),
    .CLK(clknet_leaf_20_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[45]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[45] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[1] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[45] ),
    .CLK(clknet_leaf_21_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[46]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[46] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[1] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[46] ),
    .CLK(clknet_leaf_18_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[47]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[47] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[1] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[47] ),
    .CLK(clknet_leaf_21_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[48]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[48] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[1] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[48] ),
    .CLK(clknet_leaf_31_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[49]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[49] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[1] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[49] ),
    .CLK(clknet_leaf_31_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[4]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[4] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[4] ),
    .CLK(clknet_leaf_28_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[50]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[50] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[1] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[50] ),
    .CLK(clknet_leaf_26_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[51]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[51] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[1] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[51] ),
    .CLK(clknet_leaf_26_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[52]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[52] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[1] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[52] ),
    .CLK(clknet_leaf_27_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[53]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[53] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[1] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[53] ),
    .CLK(clknet_leaf_26_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[54]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[54] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[1] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[54] ),
    .CLK(clknet_leaf_27_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[55]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[55] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[1] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[55] ),
    .CLK(clknet_leaf_24_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[56]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[56] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[1] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[56] ),
    .CLK(clknet_leaf_25_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[57]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[57] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[1] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[57] ),
    .CLK(clknet_leaf_23_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[58]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[58] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[1] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[58] ),
    .CLK(clknet_leaf_25_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[59]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[59] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[1] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[59] ),
    .CLK(clknet_leaf_23_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[5]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[5] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[5] ),
    .CLK(clknet_leaf_25_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[60]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[60] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[1] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[60] ),
    .CLK(clknet_leaf_22_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[61]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[61] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[1] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[61] ),
    .CLK(clknet_leaf_22_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[62]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[62] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[1] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[62] ),
    .CLK(clknet_leaf_23_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[63]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[63] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[1] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[63] ),
    .CLK(clknet_leaf_23_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[64]$_DFFE_PP_  (.D(net158),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[2] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[64] ),
    .CLK(clknet_leaf_29_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[65]$_DFFE_PP_  (.D(net169),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[2] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[65] ),
    .CLK(clknet_leaf_30_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[66]$_DFFE_PP_  (.D(net180),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[2] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[66] ),
    .CLK(clknet_leaf_29_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[67]$_DFFE_PP_  (.D(net183),
    .DE(net10),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[67] ),
    .CLK(clknet_leaf_27_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[68]$_DFFE_PP_  (.D(net184),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[2] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[68] ),
    .CLK(clknet_leaf_29_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[69]$_DFFE_PP_  (.D(net185),
    .DE(net9),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[69] ),
    .CLK(clknet_leaf_23_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[6]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[6] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[6] ),
    .CLK(clknet_leaf_28_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[70]$_DFFE_PP_  (.D(net186),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[2] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[70] ),
    .CLK(clknet_leaf_27_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[71]$_DFFE_PP_  (.D(net187),
    .DE(net9),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[71] ),
    .CLK(clknet_leaf_22_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[72]$_DFFE_PP_  (.D(net188),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[2] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[72] ),
    .CLK(clknet_leaf_28_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[73]$_DFFE_PP_  (.D(net189),
    .DE(net9),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[73] ),
    .CLK(clknet_leaf_21_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[74]$_DFFE_PP_  (.D(net159),
    .DE(net9),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[74] ),
    .CLK(clknet_leaf_24_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[75]$_DFFE_PP_  (.D(net160),
    .DE(net9),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[75] ),
    .CLK(clknet_leaf_24_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[76]$_DFFE_PP_  (.D(net161),
    .DE(net9),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[76] ),
    .CLK(clknet_leaf_20_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[77]$_DFFE_PP_  (.D(net162),
    .DE(net9),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[77] ),
    .CLK(clknet_leaf_21_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[78]$_DFFE_PP_  (.D(net163),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[2] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[78] ),
    .CLK(clknet_leaf_18_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[79]$_DFFE_PP_  (.D(net164),
    .DE(net9),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[79] ),
    .CLK(clknet_leaf_21_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[7]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[7] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[7] ),
    .CLK(clknet_leaf_21_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[80]$_DFFE_PP_  (.D(net165),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[2] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[80] ),
    .CLK(clknet_leaf_31_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[81]$_DFFE_PP_  (.D(net166),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[2] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[81] ),
    .CLK(clknet_leaf_31_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[82]$_DFFE_PP_  (.D(net167),
    .DE(net10),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[82] ),
    .CLK(clknet_leaf_26_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[83]$_DFFE_PP_  (.D(net168),
    .DE(net10),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[83] ),
    .CLK(clknet_leaf_26_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[84]$_DFFE_PP_  (.D(net170),
    .DE(net10),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[84] ),
    .CLK(clknet_leaf_27_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[85]$_DFFE_PP_  (.D(net171),
    .DE(net10),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[85] ),
    .CLK(clknet_leaf_26_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[86]$_DFFE_PP_  (.D(net172),
    .DE(net10),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[86] ),
    .CLK(clknet_leaf_25_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[87]$_DFFE_PP_  (.D(net173),
    .DE(net9),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[87] ),
    .CLK(clknet_leaf_23_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[88]$_DFFE_PP_  (.D(net174),
    .DE(net10),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[88] ),
    .CLK(clknet_leaf_25_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[89]$_DFFE_PP_  (.D(net175),
    .DE(net10),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[89] ),
    .CLK(clknet_leaf_23_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[8]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[8] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[8] ),
    .CLK(clknet_leaf_17_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[90]$_DFFE_PP_  (.D(net176),
    .DE(net10),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[90] ),
    .CLK(clknet_leaf_25_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[91]$_DFFE_PP_  (.D(net177),
    .DE(net10),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[91] ),
    .CLK(clknet_leaf_25_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[92]$_DFFE_PP_  (.D(net178),
    .DE(net9),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[92] ),
    .CLK(clknet_leaf_22_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[93]$_DFFE_PP_  (.D(net179),
    .DE(net9),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[93] ),
    .CLK(clknet_leaf_22_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[94]$_DFFE_PP_  (.D(net181),
    .DE(net9),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[94] ),
    .CLK(clknet_leaf_23_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[95]$_DFFE_PP_  (.D(net182),
    .DE(net9),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[95] ),
    .CLK(clknet_leaf_22_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[9]$_DFFE_PP_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_d[9] ),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[0] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.rdata_q[9] ),
    .CLK(clknet_leaf_21_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0]$_DFF_PN0_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[0] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[0] ),
    .RESET_B(net197),
    .CLK(clknet_leaf_31_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[1]$_DFF_PN0_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[1] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[0] ),
    .RESET_B(net197),
    .CLK(clknet_leaf_30_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_q[2]$_DFF_PN0_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.valid_d[2] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.fifo_busy[1] ),
    .RESET_B(net197),
    .CLK(clknet_leaf_30_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0]$_DFF_PN0_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[0] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[0] ),
    .RESET_B(net197),
    .CLK(clknet_leaf_30_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1]$_DFF_PN0_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_s[1] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.rdata_outstanding_q[1] ),
    .RESET_B(net197),
    .CLK(clknet_leaf_30_clk_i));
 sky130_fd_sc_hd__dfrtp_4 \gen_prefetch_buffer.prefetch_buffer_i.rdata_pmp_err_q[0]$_DFF_PN0_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.rdata_pmp_err_s[0] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.rdata_pmp_err_q[0] ),
    .RESET_B(net197),
    .CLK(clknet_leaf_30_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \gen_prefetch_buffer.prefetch_buffer_i.rdata_pmp_err_q[1]$_DFF_PN0_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.rdata_pmp_err_s[1] ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.rdata_pmp_err_q[1] ),
    .RESET_B(net197),
    .CLK(clknet_leaf_34_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[10]$_DFFE_PP_  (.D(net201),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[10] ),
    .CLK(clknet_leaf_33_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[11]$_DFFE_PP_  (.D(net202),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[11] ),
    .CLK(clknet_leaf_34_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[12]$_DFFE_PP_  (.D(net203),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[12] ),
    .CLK(clknet_leaf_33_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[13]$_DFFE_PP_  (.D(net204),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[13] ),
    .CLK(clknet_leaf_33_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[14]$_DFFE_PP_  (.D(net205),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[14] ),
    .CLK(clknet_leaf_32_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[15]$_DFFE_PP_  (.D(net206),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[15] ),
    .CLK(clknet_leaf_33_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[16]$_DFFE_PP_  (.D(net207),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[16] ),
    .CLK(clknet_leaf_33_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[17]$_DFFE_PP_  (.D(net208),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[17] ),
    .CLK(clknet_leaf_33_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[18]$_DFFE_PP_  (.D(net209),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[18] ),
    .CLK(clknet_leaf_32_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[19]$_DFFE_PP_  (.D(net210),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[19] ),
    .CLK(clknet_leaf_32_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[20]$_DFFE_PP_  (.D(net211),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[20] ),
    .CLK(clknet_leaf_32_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[21]$_DFFE_PP_  (.D(net212),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[21] ),
    .CLK(clknet_leaf_3_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[22]$_DFFE_PP_  (.D(net213),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[22] ),
    .CLK(clknet_leaf_32_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[23]$_DFFE_PP_  (.D(net214),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[23] ),
    .CLK(clknet_leaf_2_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[24]$_DFFE_PP_  (.D(net215),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[24] ),
    .CLK(clknet_leaf_33_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[25]$_DFFE_PP_  (.D(net216),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[25] ),
    .CLK(clknet_leaf_33_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[26]$_DFFE_PP_  (.D(net217),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[26] ),
    .CLK(clknet_leaf_32_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[27]$_DFFE_PP_  (.D(net218),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[27] ),
    .CLK(clknet_leaf_33_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[28]$_DFFE_PP_  (.D(net219),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[28] ),
    .CLK(clknet_leaf_4_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[29]$_DFFE_PP_  (.D(net220),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[29] ),
    .CLK(clknet_leaf_4_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[2]$_DFFE_PP_  (.D(net221),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[2] ),
    .CLK(clknet_leaf_0_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[30]$_DFFE_PP_  (.D(net222),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[30] ),
    .CLK(clknet_leaf_2_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[31]$_DFFE_PP_  (.D(net223),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[31] ),
    .CLK(clknet_leaf_8_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[3]$_DFFE_PP_  (.D(net224),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[3] ),
    .CLK(clknet_leaf_2_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[4]$_DFFE_PP_  (.D(net225),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[4] ),
    .CLK(clknet_leaf_0_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[5]$_DFFE_PP_  (.D(net226),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[5] ),
    .CLK(clknet_leaf_0_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[6]$_DFFE_PP_  (.D(net227),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[6] ),
    .CLK(clknet_leaf_1_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[7]$_DFFE_PP_  (.D(net228),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[7] ),
    .CLK(clknet_leaf_0_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[8]$_DFFE_PP_  (.D(net229),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[8] ),
    .CLK(clknet_leaf_0_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[9]$_DFFE_PP_  (.D(net230),
    .DE(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_en ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.stored_addr_q[9] ),
    .CLK(clknet_leaf_0_clk_i));
 sky130_fd_sc_hd__dfrtp_1 \gen_prefetch_buffer.prefetch_buffer_i.valid_req_q$_DFF_PN0_  (.D(\gen_prefetch_buffer.prefetch_buffer_i.valid_req_d ),
    .Q(\gen_prefetch_buffer.prefetch_buffer_i.valid_req_q ),
    .RESET_B(net197),
    .CLK(clknet_leaf_34_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \illegal_c_insn_id_o$_DFFE_PP_  (.D(\compressed_decoder_i.illegal_instr_o ),
    .DE(net7),
    .Q(net200),
    .CLK(clknet_leaf_14_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_fetch_err_o$_DFFE_PP_  (.D(fetch_err),
    .DE(net7),
    .Q(net231),
    .CLK(clknet_leaf_29_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_fetch_err_plus2_o$_SDFFCE_PN0P_  (.D(_0000_),
    .DE(net7),
    .Q(net232),
    .CLK(clknet_leaf_29_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_is_compressed_id_o$_DFFE_PP_  (.D(\compressed_decoder_i.is_compressed_o ),
    .DE(net6),
    .Q(net233),
    .CLK(clknet_leaf_19_clk_i));
 sky130_fd_sc_hd__dfrtp_2 \instr_new_id_q$_DFF_PN0_  (.D(net7),
    .Q(net234),
    .RESET_B(net197),
    .CLK(clknet_leaf_29_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_rdata_alu_id_o[0]$_DFFE_PP_  (.D(\compressed_decoder_i.instr_o[0] ),
    .DE(net6),
    .Q(net235),
    .CLK(clknet_leaf_19_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_rdata_alu_id_o[10]$_DFFE_PP_  (.D(\compressed_decoder_i.instr_o[10] ),
    .DE(net7),
    .Q(net236),
    .CLK(clknet_leaf_14_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_rdata_alu_id_o[11]$_DFFE_PP_  (.D(\compressed_decoder_i.instr_o[11] ),
    .DE(net6),
    .Q(net237),
    .CLK(clknet_leaf_14_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_rdata_alu_id_o[12]$_DFFE_PP_  (.D(\compressed_decoder_i.instr_o[12] ),
    .DE(net6),
    .Q(net238),
    .CLK(clknet_leaf_14_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_rdata_alu_id_o[13]$_DFFE_PP_  (.D(\compressed_decoder_i.instr_o[13] ),
    .DE(net6),
    .Q(net239),
    .CLK(clknet_leaf_13_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_rdata_alu_id_o[14]$_DFFE_PP_  (.D(\compressed_decoder_i.instr_o[14] ),
    .DE(net6),
    .Q(net240),
    .CLK(clknet_leaf_14_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_rdata_alu_id_o[15]$_DFFE_PP_  (.D(\compressed_decoder_i.instr_o[15] ),
    .DE(net6),
    .Q(net241),
    .CLK(clknet_leaf_15_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_rdata_alu_id_o[16]$_DFFE_PP_  (.D(\compressed_decoder_i.instr_o[16] ),
    .DE(net6),
    .Q(net242),
    .CLK(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_rdata_alu_id_o[17]$_DFFE_PP_  (.D(\compressed_decoder_i.instr_o[17] ),
    .DE(net6),
    .Q(net243),
    .CLK(clknet_leaf_17_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_rdata_alu_id_o[18]$_DFFE_PP_  (.D(\compressed_decoder_i.instr_o[18] ),
    .DE(net6),
    .Q(net244),
    .CLK(clknet_leaf_19_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_rdata_alu_id_o[19]$_DFFE_PP_  (.D(\compressed_decoder_i.instr_o[19] ),
    .DE(net6),
    .Q(net245),
    .CLK(clknet_leaf_19_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_rdata_alu_id_o[1]$_DFFE_PP_  (.D(\compressed_decoder_i.instr_o[1] ),
    .DE(net7),
    .Q(net246),
    .CLK(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_rdata_alu_id_o[20]$_DFFE_PP_  (.D(\compressed_decoder_i.instr_o[20] ),
    .DE(net7),
    .Q(net247),
    .CLK(clknet_leaf_17_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_rdata_alu_id_o[21]$_DFFE_PP_  (.D(\compressed_decoder_i.instr_o[21] ),
    .DE(net6),
    .Q(net248),
    .CLK(clknet_leaf_16_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_rdata_alu_id_o[22]$_DFFE_PP_  (.D(\compressed_decoder_i.instr_o[22] ),
    .DE(net6),
    .Q(net249),
    .CLK(clknet_leaf_15_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_rdata_alu_id_o[23]$_DFFE_PP_  (.D(\compressed_decoder_i.instr_o[23] ),
    .DE(net6),
    .Q(net250),
    .CLK(clknet_leaf_16_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_rdata_alu_id_o[24]$_DFFE_PP_  (.D(\compressed_decoder_i.instr_o[24] ),
    .DE(net6),
    .Q(net251),
    .CLK(clknet_leaf_15_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_rdata_alu_id_o[25]$_DFFE_PP_  (.D(\compressed_decoder_i.instr_o[25] ),
    .DE(net6),
    .Q(net252),
    .CLK(clknet_leaf_19_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_rdata_alu_id_o[26]$_DFFE_PP_  (.D(\compressed_decoder_i.instr_o[26] ),
    .DE(net6),
    .Q(net253),
    .CLK(clknet_leaf_19_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_rdata_alu_id_o[27]$_DFFE_PP_  (.D(\compressed_decoder_i.instr_o[27] ),
    .DE(net6),
    .Q(net254),
    .CLK(clknet_leaf_20_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_rdata_alu_id_o[28]$_DFFE_PP_  (.D(\compressed_decoder_i.instr_o[28] ),
    .DE(net6),
    .Q(net255),
    .CLK(clknet_leaf_20_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_rdata_alu_id_o[29]$_DFFE_PP_  (.D(\compressed_decoder_i.instr_o[29] ),
    .DE(net6),
    .Q(net256),
    .CLK(clknet_leaf_19_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_rdata_alu_id_o[2]$_DFFE_PP_  (.D(\compressed_decoder_i.instr_o[2] ),
    .DE(net7),
    .Q(net257),
    .CLK(clknet_leaf_14_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_rdata_alu_id_o[30]$_DFFE_PP_  (.D(\compressed_decoder_i.instr_o[30] ),
    .DE(net6),
    .Q(net258),
    .CLK(clknet_leaf_19_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_rdata_alu_id_o[31]$_DFFE_PP_  (.D(\compressed_decoder_i.instr_o[31] ),
    .DE(net6),
    .Q(net259),
    .CLK(clknet_leaf_15_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_rdata_alu_id_o[3]$_DFFE_PP_  (.D(\compressed_decoder_i.instr_o[3] ),
    .DE(net6),
    .Q(net260),
    .CLK(clknet_leaf_15_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_rdata_alu_id_o[4]$_DFFE_PP_  (.D(\compressed_decoder_i.instr_o[4] ),
    .DE(net6),
    .Q(net261),
    .CLK(clknet_leaf_13_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_rdata_alu_id_o[5]$_DFFE_PP_  (.D(\compressed_decoder_i.instr_o[5] ),
    .DE(net6),
    .Q(net262),
    .CLK(clknet_leaf_15_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_rdata_alu_id_o[6]$_DFFE_PP_  (.D(\compressed_decoder_i.instr_o[6] ),
    .DE(net6),
    .Q(net263),
    .CLK(clknet_leaf_15_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_rdata_alu_id_o[7]$_DFFE_PP_  (.D(\compressed_decoder_i.instr_o[7] ),
    .DE(net6),
    .Q(net264),
    .CLK(clknet_leaf_13_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_rdata_alu_id_o[8]$_DFFE_PP_  (.D(\compressed_decoder_i.instr_o[8] ),
    .DE(net7),
    .Q(net265),
    .CLK(clknet_leaf_13_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_rdata_alu_id_o[9]$_DFFE_PP_  (.D(\compressed_decoder_i.instr_o[9] ),
    .DE(net6),
    .Q(net266),
    .CLK(clknet_leaf_13_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_rdata_c_id_o[0]$_DFFE_PP_  (.D(\compressed_decoder_i.instr_i[0] ),
    .DE(net6),
    .Q(net267),
    .CLK(clknet_leaf_13_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_rdata_c_id_o[10]$_DFFE_PP_  (.D(\compressed_decoder_i.instr_i[10] ),
    .DE(net6),
    .Q(net268),
    .CLK(clknet_leaf_20_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_rdata_c_id_o[11]$_DFFE_PP_  (.D(\compressed_decoder_i.instr_i[11] ),
    .DE(net6),
    .Q(net269),
    .CLK(clknet_leaf_20_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_rdata_c_id_o[12]$_DFFE_PP_  (.D(\compressed_decoder_i.instr_i[12] ),
    .DE(net6),
    .Q(net270),
    .CLK(clknet_leaf_19_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_rdata_c_id_o[13]$_DFFE_PP_  (.D(\compressed_decoder_i.instr_i[13] ),
    .DE(net6),
    .Q(net271),
    .CLK(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_rdata_c_id_o[14]$_DFFE_PP_  (.D(\compressed_decoder_i.instr_i[14] ),
    .DE(net6),
    .Q(net272),
    .CLK(clknet_leaf_15_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_rdata_c_id_o[15]$_DFFE_PP_  (.D(\compressed_decoder_i.instr_i[15] ),
    .DE(net6),
    .Q(net273),
    .CLK(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_rdata_c_id_o[1]$_DFFE_PP_  (.D(\compressed_decoder_i.instr_i[1] ),
    .DE(net6),
    .Q(net274),
    .CLK(clknet_leaf_14_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_rdata_c_id_o[2]$_DFFE_PP_  (.D(\compressed_decoder_i.instr_i[2] ),
    .DE(net6),
    .Q(net275),
    .CLK(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_rdata_c_id_o[3]$_DFFE_PP_  (.D(\compressed_decoder_i.instr_i[3] ),
    .DE(net6),
    .Q(net276),
    .CLK(clknet_leaf_17_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_rdata_c_id_o[4]$_DFFE_PP_  (.D(\compressed_decoder_i.instr_i[4] ),
    .DE(net6),
    .Q(net277),
    .CLK(clknet_leaf_17_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_rdata_c_id_o[5]$_DFFE_PP_  (.D(\compressed_decoder_i.instr_i[5] ),
    .DE(net6),
    .Q(net278),
    .CLK(clknet_leaf_14_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_rdata_c_id_o[6]$_DFFE_PP_  (.D(\compressed_decoder_i.instr_i[6] ),
    .DE(net6),
    .Q(net279),
    .CLK(clknet_leaf_14_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_rdata_c_id_o[7]$_DFFE_PP_  (.D(\compressed_decoder_i.instr_i[7] ),
    .DE(net6),
    .Q(net280),
    .CLK(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_rdata_c_id_o[8]$_DFFE_PP_  (.D(\compressed_decoder_i.instr_i[8] ),
    .DE(net7),
    .Q(net281),
    .CLK(clknet_leaf_16_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \instr_rdata_c_id_o[9]$_DFFE_PP_  (.D(\compressed_decoder_i.instr_i[9] ),
    .DE(net6),
    .Q(net282),
    .CLK(clknet_leaf_18_clk_i));
 sky130_fd_sc_hd__dfrtp_2 \instr_valid_id_q$_DFF_PN0_  (.D(instr_valid_id_d),
    .Q(net316),
    .RESET_B(net197),
    .CLK(clknet_leaf_0_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \pc_id_o[10]$_DFFE_PP_  (.D(net348),
    .DE(net7),
    .Q(net317),
    .CLK(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \pc_id_o[11]$_DFFE_PP_  (.D(net349),
    .DE(net7),
    .Q(net318),
    .CLK(clknet_leaf_11_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \pc_id_o[12]$_DFFE_PP_  (.D(net350),
    .DE(net7),
    .Q(net319),
    .CLK(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \pc_id_o[13]$_DFFE_PP_  (.D(net351),
    .DE(net7),
    .Q(net320),
    .CLK(clknet_leaf_11_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \pc_id_o[14]$_DFFE_PP_  (.D(net352),
    .DE(net7),
    .Q(net321),
    .CLK(clknet_leaf_9_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \pc_id_o[15]$_DFFE_PP_  (.D(net353),
    .DE(net7),
    .Q(net322),
    .CLK(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \pc_id_o[16]$_DFFE_PP_  (.D(net354),
    .DE(net7),
    .Q(net323),
    .CLK(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \pc_id_o[17]$_DFFE_PP_  (.D(net355),
    .DE(net7),
    .Q(net324),
    .CLK(clknet_leaf_7_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \pc_id_o[18]$_DFFE_PP_  (.D(net356),
    .DE(if_id_pipe_reg_we),
    .Q(net325),
    .CLK(clknet_leaf_5_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \pc_id_o[19]$_DFFE_PP_  (.D(net357),
    .DE(if_id_pipe_reg_we),
    .Q(net326),
    .CLK(clknet_leaf_5_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \pc_id_o[1]$_DFFE_PP_  (.D(net358),
    .DE(net7),
    .Q(net327),
    .CLK(clknet_leaf_29_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \pc_id_o[20]$_DFFE_PP_  (.D(net359),
    .DE(if_id_pipe_reg_we),
    .Q(net328),
    .CLK(clknet_leaf_5_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \pc_id_o[21]$_DFFE_PP_  (.D(net360),
    .DE(if_id_pipe_reg_we),
    .Q(net329),
    .CLK(clknet_leaf_5_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \pc_id_o[22]$_DFFE_PP_  (.D(net361),
    .DE(net7),
    .Q(net330),
    .CLK(clknet_leaf_11_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \pc_id_o[23]$_DFFE_PP_  (.D(net362),
    .DE(net7),
    .Q(net331),
    .CLK(clknet_leaf_12_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \pc_id_o[24]$_DFFE_PP_  (.D(net363),
    .DE(net7),
    .Q(net332),
    .CLK(clknet_leaf_12_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \pc_id_o[25]$_DFFE_PP_  (.D(net364),
    .DE(net7),
    .Q(net333),
    .CLK(clknet_leaf_12_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \pc_id_o[26]$_DFFE_PP_  (.D(net365),
    .DE(net7),
    .Q(net334),
    .CLK(clknet_leaf_12_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \pc_id_o[27]$_DFFE_PP_  (.D(net366),
    .DE(net7),
    .Q(net335),
    .CLK(clknet_leaf_12_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \pc_id_o[28]$_DFFE_PP_  (.D(net367),
    .DE(net7),
    .Q(net336),
    .CLK(clknet_leaf_6_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \pc_id_o[29]$_DFFE_PP_  (.D(net368),
    .DE(net7),
    .Q(net337),
    .CLK(clknet_leaf_6_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \pc_id_o[2]$_DFFE_PP_  (.D(net369),
    .DE(net7),
    .Q(net338),
    .CLK(clknet_leaf_17_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \pc_id_o[30]$_DFFE_PP_  (.D(net370),
    .DE(net7),
    .Q(net339),
    .CLK(clknet_leaf_6_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \pc_id_o[31]$_DFFE_PP_  (.D(net371),
    .DE(if_id_pipe_reg_we),
    .Q(net340),
    .CLK(clknet_leaf_5_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \pc_id_o[3]$_DFFE_PP_  (.D(net372),
    .DE(net7),
    .Q(net341),
    .CLK(clknet_leaf_9_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \pc_id_o[4]$_DFFE_PP_  (.D(net373),
    .DE(net7),
    .Q(net342),
    .CLK(clknet_leaf_16_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \pc_id_o[5]$_DFFE_PP_  (.D(net374),
    .DE(net6),
    .Q(net343),
    .CLK(clknet_leaf_16_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \pc_id_o[6]$_DFFE_PP_  (.D(net375),
    .DE(net6),
    .Q(net344),
    .CLK(clknet_leaf_9_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \pc_id_o[7]$_DFFE_PP_  (.D(net376),
    .DE(net6),
    .Q(net345),
    .CLK(clknet_leaf_16_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \pc_id_o[8]$_DFFE_PP_  (.D(net377),
    .DE(net7),
    .Q(net346),
    .CLK(clknet_leaf_9_clk_i));
 sky130_fd_sc_hd__edfxtp_1 \pc_id_o[9]$_DFFE_PP_  (.D(net378),
    .DE(net7),
    .Q(net347),
    .CLK(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1143 ();
 sky130_fd_sc_hd__buf_16 load_slew6 (.A(net7),
    .X(net6));
 sky130_fd_sc_hd__buf_12 load_slew7 (.A(if_id_pipe_reg_we),
    .X(net7));
 sky130_fd_sc_hd__buf_2 wire8 (.A(_1053_),
    .X(net8));
 sky130_fd_sc_hd__buf_6 wire9 (.A(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[2] ),
    .X(net9));
 sky130_fd_sc_hd__buf_6 load_slew10 (.A(\gen_prefetch_buffer.prefetch_buffer_i.fifo_i.entry_en[2] ),
    .X(net10));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input1 (.A(boot_addr_i[10]),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input2 (.A(boot_addr_i[11]),
    .X(net2));
 sky130_fd_sc_hd__buf_2 input3 (.A(boot_addr_i[12]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input4 (.A(boot_addr_i[13]),
    .X(net4));
 sky130_fd_sc_hd__buf_4 input5 (.A(boot_addr_i[14]),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input6 (.A(boot_addr_i[15]),
    .X(net11));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input7 (.A(boot_addr_i[16]),
    .X(net12));
 sky130_fd_sc_hd__buf_4 input8 (.A(boot_addr_i[17]),
    .X(net13));
 sky130_fd_sc_hd__buf_4 input9 (.A(boot_addr_i[18]),
    .X(net14));
 sky130_fd_sc_hd__buf_2 input10 (.A(boot_addr_i[19]),
    .X(net15));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input11 (.A(boot_addr_i[20]),
    .X(net16));
 sky130_fd_sc_hd__buf_1 input12 (.A(boot_addr_i[21]),
    .X(net17));
 sky130_fd_sc_hd__buf_1 input13 (.A(boot_addr_i[22]),
    .X(net18));
 sky130_fd_sc_hd__buf_2 input14 (.A(boot_addr_i[23]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input15 (.A(boot_addr_i[24]),
    .X(net20));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input16 (.A(boot_addr_i[25]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input17 (.A(boot_addr_i[26]),
    .X(net22));
 sky130_fd_sc_hd__buf_1 input18 (.A(boot_addr_i[27]),
    .X(net23));
 sky130_fd_sc_hd__buf_1 input19 (.A(boot_addr_i[28]),
    .X(net24));
 sky130_fd_sc_hd__buf_1 input20 (.A(boot_addr_i[29]),
    .X(net25));
 sky130_fd_sc_hd__buf_2 input21 (.A(boot_addr_i[30]),
    .X(net26));
 sky130_fd_sc_hd__buf_4 input22 (.A(boot_addr_i[31]),
    .X(net27));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input23 (.A(boot_addr_i[8]),
    .X(net28));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input24 (.A(boot_addr_i[9]),
    .X(net29));
 sky130_fd_sc_hd__buf_1 input25 (.A(branch_target_ex_i[10]),
    .X(net30));
 sky130_fd_sc_hd__buf_1 input26 (.A(branch_target_ex_i[11]),
    .X(net31));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input27 (.A(branch_target_ex_i[12]),
    .X(net32));
 sky130_fd_sc_hd__buf_1 input28 (.A(branch_target_ex_i[13]),
    .X(net33));
 sky130_fd_sc_hd__buf_2 input29 (.A(branch_target_ex_i[14]),
    .X(net34));
 sky130_fd_sc_hd__buf_2 input30 (.A(branch_target_ex_i[15]),
    .X(net35));
 sky130_fd_sc_hd__buf_2 input31 (.A(branch_target_ex_i[16]),
    .X(net36));
 sky130_fd_sc_hd__buf_2 input32 (.A(branch_target_ex_i[17]),
    .X(net37));
 sky130_fd_sc_hd__buf_1 input33 (.A(branch_target_ex_i[18]),
    .X(net38));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input34 (.A(branch_target_ex_i[19]),
    .X(net39));
 sky130_fd_sc_hd__buf_2 input35 (.A(branch_target_ex_i[1]),
    .X(net40));
 sky130_fd_sc_hd__buf_1 input36 (.A(branch_target_ex_i[20]),
    .X(net41));
 sky130_fd_sc_hd__buf_1 input37 (.A(branch_target_ex_i[21]),
    .X(net42));
 sky130_fd_sc_hd__buf_1 input38 (.A(branch_target_ex_i[22]),
    .X(net43));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input39 (.A(branch_target_ex_i[23]),
    .X(net44));
 sky130_fd_sc_hd__buf_1 input40 (.A(branch_target_ex_i[24]),
    .X(net45));
 sky130_fd_sc_hd__buf_1 input41 (.A(branch_target_ex_i[25]),
    .X(net46));
 sky130_fd_sc_hd__buf_2 input42 (.A(branch_target_ex_i[26]),
    .X(net47));
 sky130_fd_sc_hd__buf_1 input43 (.A(branch_target_ex_i[27]),
    .X(net48));
 sky130_fd_sc_hd__buf_1 input44 (.A(branch_target_ex_i[28]),
    .X(net49));
 sky130_fd_sc_hd__buf_1 input45 (.A(branch_target_ex_i[29]),
    .X(net50));
 sky130_fd_sc_hd__buf_1 input46 (.A(branch_target_ex_i[2]),
    .X(net51));
 sky130_fd_sc_hd__buf_2 input47 (.A(branch_target_ex_i[30]),
    .X(net52));
 sky130_fd_sc_hd__buf_4 input48 (.A(branch_target_ex_i[31]),
    .X(net53));
 sky130_fd_sc_hd__buf_1 input49 (.A(branch_target_ex_i[3]),
    .X(net54));
 sky130_fd_sc_hd__buf_2 input50 (.A(branch_target_ex_i[4]),
    .X(net55));
 sky130_fd_sc_hd__buf_2 input51 (.A(branch_target_ex_i[5]),
    .X(net56));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input52 (.A(branch_target_ex_i[6]),
    .X(net57));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input53 (.A(branch_target_ex_i[7]),
    .X(net58));
 sky130_fd_sc_hd__buf_1 input54 (.A(branch_target_ex_i[8]),
    .X(net59));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input55 (.A(branch_target_ex_i[9]),
    .X(net60));
 sky130_fd_sc_hd__buf_1 input56 (.A(csr_depc_i[10]),
    .X(net61));
 sky130_fd_sc_hd__buf_1 input57 (.A(csr_depc_i[11]),
    .X(net62));
 sky130_fd_sc_hd__buf_1 input58 (.A(csr_depc_i[12]),
    .X(net63));
 sky130_fd_sc_hd__buf_1 input59 (.A(csr_depc_i[13]),
    .X(net64));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input60 (.A(csr_depc_i[14]),
    .X(net65));
 sky130_fd_sc_hd__buf_1 input61 (.A(csr_depc_i[15]),
    .X(net66));
 sky130_fd_sc_hd__buf_1 input62 (.A(csr_depc_i[16]),
    .X(net67));
 sky130_fd_sc_hd__buf_4 input63 (.A(csr_depc_i[17]),
    .X(net68));
 sky130_fd_sc_hd__buf_4 input64 (.A(csr_depc_i[18]),
    .X(net69));
 sky130_fd_sc_hd__buf_2 input65 (.A(csr_depc_i[19]),
    .X(net70));
 sky130_fd_sc_hd__buf_2 input66 (.A(csr_depc_i[1]),
    .X(net71));
 sky130_fd_sc_hd__buf_1 input67 (.A(csr_depc_i[20]),
    .X(net72));
 sky130_fd_sc_hd__buf_1 input68 (.A(csr_depc_i[21]),
    .X(net73));
 sky130_fd_sc_hd__buf_1 input69 (.A(csr_depc_i[22]),
    .X(net74));
 sky130_fd_sc_hd__buf_2 input70 (.A(csr_depc_i[23]),
    .X(net75));
 sky130_fd_sc_hd__buf_1 input71 (.A(csr_depc_i[24]),
    .X(net76));
 sky130_fd_sc_hd__buf_1 input72 (.A(csr_depc_i[25]),
    .X(net77));
 sky130_fd_sc_hd__buf_4 input73 (.A(csr_depc_i[26]),
    .X(net78));
 sky130_fd_sc_hd__buf_1 input74 (.A(csr_depc_i[27]),
    .X(net79));
 sky130_fd_sc_hd__buf_1 input75 (.A(csr_depc_i[28]),
    .X(net80));
 sky130_fd_sc_hd__buf_1 input76 (.A(csr_depc_i[29]),
    .X(net81));
 sky130_fd_sc_hd__buf_2 input77 (.A(csr_depc_i[2]),
    .X(net82));
 sky130_fd_sc_hd__buf_1 input78 (.A(csr_depc_i[30]),
    .X(net83));
 sky130_fd_sc_hd__buf_2 input79 (.A(csr_depc_i[31]),
    .X(net84));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input80 (.A(csr_depc_i[3]),
    .X(net85));
 sky130_fd_sc_hd__buf_4 input81 (.A(csr_depc_i[4]),
    .X(net86));
 sky130_fd_sc_hd__buf_2 input82 (.A(csr_depc_i[5]),
    .X(net87));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input83 (.A(csr_depc_i[6]),
    .X(net88));
 sky130_fd_sc_hd__buf_1 input84 (.A(csr_depc_i[7]),
    .X(net89));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input85 (.A(csr_depc_i[8]),
    .X(net90));
 sky130_fd_sc_hd__buf_1 input86 (.A(csr_depc_i[9]),
    .X(net91));
 sky130_fd_sc_hd__buf_1 input87 (.A(csr_mepc_i[10]),
    .X(net92));
 sky130_fd_sc_hd__buf_1 input88 (.A(csr_mepc_i[11]),
    .X(net93));
 sky130_fd_sc_hd__buf_2 input89 (.A(csr_mepc_i[12]),
    .X(net94));
 sky130_fd_sc_hd__buf_1 input90 (.A(csr_mepc_i[13]),
    .X(net95));
 sky130_fd_sc_hd__buf_2 input91 (.A(csr_mepc_i[14]),
    .X(net96));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input92 (.A(csr_mepc_i[15]),
    .X(net97));
 sky130_fd_sc_hd__buf_1 input93 (.A(csr_mepc_i[16]),
    .X(net98));
 sky130_fd_sc_hd__buf_2 input94 (.A(csr_mepc_i[17]),
    .X(net99));
 sky130_fd_sc_hd__buf_1 input95 (.A(csr_mepc_i[18]),
    .X(net100));
 sky130_fd_sc_hd__buf_2 input96 (.A(csr_mepc_i[19]),
    .X(net101));
 sky130_fd_sc_hd__buf_2 input97 (.A(csr_mepc_i[1]),
    .X(net102));
 sky130_fd_sc_hd__buf_2 input98 (.A(csr_mepc_i[20]),
    .X(net103));
 sky130_fd_sc_hd__buf_1 input99 (.A(csr_mepc_i[21]),
    .X(net104));
 sky130_fd_sc_hd__buf_1 input100 (.A(csr_mepc_i[22]),
    .X(net105));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input101 (.A(csr_mepc_i[23]),
    .X(net106));
 sky130_fd_sc_hd__buf_1 input102 (.A(csr_mepc_i[24]),
    .X(net107));
 sky130_fd_sc_hd__buf_1 input103 (.A(csr_mepc_i[25]),
    .X(net108));
 sky130_fd_sc_hd__buf_1 input104 (.A(csr_mepc_i[26]),
    .X(net109));
 sky130_fd_sc_hd__buf_1 input105 (.A(csr_mepc_i[27]),
    .X(net110));
 sky130_fd_sc_hd__buf_1 input106 (.A(csr_mepc_i[28]),
    .X(net111));
 sky130_fd_sc_hd__buf_1 input107 (.A(csr_mepc_i[29]),
    .X(net112));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input108 (.A(csr_mepc_i[2]),
    .X(net113));
 sky130_fd_sc_hd__buf_1 input109 (.A(csr_mepc_i[30]),
    .X(net114));
 sky130_fd_sc_hd__buf_4 input110 (.A(csr_mepc_i[31]),
    .X(net115));
 sky130_fd_sc_hd__buf_2 input111 (.A(csr_mepc_i[3]),
    .X(net116));
 sky130_fd_sc_hd__buf_2 input112 (.A(csr_mepc_i[4]),
    .X(net117));
 sky130_fd_sc_hd__buf_1 input113 (.A(csr_mepc_i[5]),
    .X(net118));
 sky130_fd_sc_hd__buf_2 input114 (.A(csr_mepc_i[6]),
    .X(net119));
 sky130_fd_sc_hd__buf_1 input115 (.A(csr_mepc_i[7]),
    .X(net120));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input116 (.A(csr_mepc_i[8]),
    .X(net121));
 sky130_fd_sc_hd__buf_1 input117 (.A(csr_mepc_i[9]),
    .X(net122));
 sky130_fd_sc_hd__buf_1 input118 (.A(csr_mtvec_i[10]),
    .X(net123));
 sky130_fd_sc_hd__buf_1 input119 (.A(csr_mtvec_i[11]),
    .X(net124));
 sky130_fd_sc_hd__buf_1 input120 (.A(csr_mtvec_i[12]),
    .X(net125));
 sky130_fd_sc_hd__buf_1 input121 (.A(csr_mtvec_i[13]),
    .X(net126));
 sky130_fd_sc_hd__buf_2 input122 (.A(csr_mtvec_i[14]),
    .X(net127));
 sky130_fd_sc_hd__buf_1 input123 (.A(csr_mtvec_i[15]),
    .X(net128));
 sky130_fd_sc_hd__buf_1 input124 (.A(csr_mtvec_i[16]),
    .X(net129));
 sky130_fd_sc_hd__buf_2 input125 (.A(csr_mtvec_i[17]),
    .X(net130));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input126 (.A(csr_mtvec_i[18]),
    .X(net131));
 sky130_fd_sc_hd__buf_2 input127 (.A(csr_mtvec_i[19]),
    .X(net132));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input128 (.A(csr_mtvec_i[20]),
    .X(net133));
 sky130_fd_sc_hd__buf_1 input129 (.A(csr_mtvec_i[21]),
    .X(net134));
 sky130_fd_sc_hd__buf_1 input130 (.A(csr_mtvec_i[22]),
    .X(net135));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input131 (.A(csr_mtvec_i[23]),
    .X(net136));
 sky130_fd_sc_hd__buf_4 input132 (.A(csr_mtvec_i[24]),
    .X(net137));
 sky130_fd_sc_hd__buf_2 input133 (.A(csr_mtvec_i[25]),
    .X(net138));
 sky130_fd_sc_hd__buf_1 input134 (.A(csr_mtvec_i[26]),
    .X(net139));
 sky130_fd_sc_hd__buf_1 input135 (.A(csr_mtvec_i[27]),
    .X(net140));
 sky130_fd_sc_hd__buf_1 input136 (.A(csr_mtvec_i[28]),
    .X(net141));
 sky130_fd_sc_hd__buf_1 input137 (.A(csr_mtvec_i[29]),
    .X(net142));
 sky130_fd_sc_hd__buf_2 input138 (.A(csr_mtvec_i[30]),
    .X(net143));
 sky130_fd_sc_hd__buf_1 input139 (.A(csr_mtvec_i[31]),
    .X(net144));
 sky130_fd_sc_hd__buf_2 input140 (.A(csr_mtvec_i[8]),
    .X(net145));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input141 (.A(csr_mtvec_i[9]),
    .X(net146));
 sky130_fd_sc_hd__buf_2 input142 (.A(exc_cause[0]),
    .X(net147));
 sky130_fd_sc_hd__buf_1 input143 (.A(exc_cause[1]),
    .X(net148));
 sky130_fd_sc_hd__buf_2 input144 (.A(exc_cause[2]),
    .X(net149));
 sky130_fd_sc_hd__buf_4 input145 (.A(exc_cause[3]),
    .X(net150));
 sky130_fd_sc_hd__buf_2 input146 (.A(exc_cause[4]),
    .X(net151));
 sky130_fd_sc_hd__buf_4 input147 (.A(exc_pc_mux_i[0]),
    .X(net152));
 sky130_fd_sc_hd__buf_2 input148 (.A(exc_pc_mux_i[1]),
    .X(net153));
 sky130_fd_sc_hd__buf_2 input149 (.A(id_in_ready_i),
    .X(net154));
 sky130_fd_sc_hd__buf_1 input150 (.A(instr_err_i),
    .X(net155));
 sky130_fd_sc_hd__buf_1 input151 (.A(instr_gnt_i),
    .X(net156));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input152 (.A(instr_pmp_err_i),
    .X(net157));
 sky130_fd_sc_hd__buf_2 input153 (.A(instr_rdata_i[0]),
    .X(net158));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input154 (.A(instr_rdata_i[10]),
    .X(net159));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input155 (.A(instr_rdata_i[11]),
    .X(net160));
 sky130_fd_sc_hd__buf_1 input156 (.A(instr_rdata_i[12]),
    .X(net161));
 sky130_fd_sc_hd__buf_1 input157 (.A(instr_rdata_i[13]),
    .X(net162));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input158 (.A(instr_rdata_i[14]),
    .X(net163));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input159 (.A(instr_rdata_i[15]),
    .X(net164));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input160 (.A(instr_rdata_i[16]),
    .X(net165));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input161 (.A(instr_rdata_i[17]),
    .X(net166));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input162 (.A(instr_rdata_i[18]),
    .X(net167));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input163 (.A(instr_rdata_i[19]),
    .X(net168));
 sky130_fd_sc_hd__buf_2 input164 (.A(instr_rdata_i[1]),
    .X(net169));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input165 (.A(instr_rdata_i[20]),
    .X(net170));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input166 (.A(instr_rdata_i[21]),
    .X(net171));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input167 (.A(instr_rdata_i[22]),
    .X(net172));
 sky130_fd_sc_hd__buf_1 input168 (.A(instr_rdata_i[23]),
    .X(net173));
 sky130_fd_sc_hd__buf_1 input169 (.A(instr_rdata_i[24]),
    .X(net174));
 sky130_fd_sc_hd__buf_1 input170 (.A(instr_rdata_i[25]),
    .X(net175));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input171 (.A(instr_rdata_i[26]),
    .X(net176));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input172 (.A(instr_rdata_i[27]),
    .X(net177));
 sky130_fd_sc_hd__buf_1 input173 (.A(instr_rdata_i[28]),
    .X(net178));
 sky130_fd_sc_hd__buf_1 input174 (.A(instr_rdata_i[29]),
    .X(net179));
 sky130_fd_sc_hd__buf_2 input175 (.A(instr_rdata_i[2]),
    .X(net180));
 sky130_fd_sc_hd__buf_1 input176 (.A(instr_rdata_i[30]),
    .X(net181));
 sky130_fd_sc_hd__buf_1 input177 (.A(instr_rdata_i[31]),
    .X(net182));
 sky130_fd_sc_hd__buf_1 input178 (.A(instr_rdata_i[3]),
    .X(net183));
 sky130_fd_sc_hd__clkdlybuf4s15_2 input179 (.A(instr_rdata_i[4]),
    .X(net184));
 sky130_fd_sc_hd__buf_1 input180 (.A(instr_rdata_i[5]),
    .X(net185));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input181 (.A(instr_rdata_i[6]),
    .X(net186));
 sky130_fd_sc_hd__buf_2 input182 (.A(instr_rdata_i[7]),
    .X(net187));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input183 (.A(instr_rdata_i[8]),
    .X(net188));
 sky130_fd_sc_hd__buf_1 input184 (.A(instr_rdata_i[9]),
    .X(net189));
 sky130_fd_sc_hd__buf_2 input185 (.A(instr_rvalid_i),
    .X(net190));
 sky130_fd_sc_hd__clkdlybuf4s18_2 input186 (.A(instr_valid_clear_i),
    .X(net191));
 sky130_fd_sc_hd__buf_4 input187 (.A(nt_branch_mispredict_i),
    .X(net192));
 sky130_fd_sc_hd__buf_2 input188 (.A(pc_mux_i[0]),
    .X(net193));
 sky130_fd_sc_hd__buf_2 input189 (.A(pc_mux_i[2]),
    .X(net194));
 sky130_fd_sc_hd__buf_4 input190 (.A(pc_set_i),
    .X(net195));
 sky130_fd_sc_hd__buf_1 input191 (.A(req_i),
    .X(net196));
 sky130_fd_sc_hd__buf_6 input192 (.A(rst_ni),
    .X(net197));
 sky130_fd_sc_hd__buf_1 output193 (.A(net198),
    .X(csr_mtvec_init_o));
 sky130_fd_sc_hd__buf_1 output194 (.A(net199),
    .X(if_busy_o));
 sky130_fd_sc_hd__buf_1 output195 (.A(net200),
    .X(illegal_c_insn_id_o));
 sky130_fd_sc_hd__buf_1 output196 (.A(net201),
    .X(instr_addr_o[10]));
 sky130_fd_sc_hd__buf_1 output197 (.A(net202),
    .X(instr_addr_o[11]));
 sky130_fd_sc_hd__buf_1 output198 (.A(net203),
    .X(instr_addr_o[12]));
 sky130_fd_sc_hd__buf_1 output199 (.A(net204),
    .X(instr_addr_o[13]));
 sky130_fd_sc_hd__buf_1 output200 (.A(net205),
    .X(instr_addr_o[14]));
 sky130_fd_sc_hd__buf_1 output201 (.A(net206),
    .X(instr_addr_o[15]));
 sky130_fd_sc_hd__buf_1 output202 (.A(net207),
    .X(instr_addr_o[16]));
 sky130_fd_sc_hd__buf_1 output203 (.A(net208),
    .X(instr_addr_o[17]));
 sky130_fd_sc_hd__buf_1 output204 (.A(net209),
    .X(instr_addr_o[18]));
 sky130_fd_sc_hd__buf_1 output205 (.A(net210),
    .X(instr_addr_o[19]));
 sky130_fd_sc_hd__buf_1 output206 (.A(net211),
    .X(instr_addr_o[20]));
 sky130_fd_sc_hd__buf_1 output207 (.A(net212),
    .X(instr_addr_o[21]));
 sky130_fd_sc_hd__buf_1 output208 (.A(net213),
    .X(instr_addr_o[22]));
 sky130_fd_sc_hd__buf_1 output209 (.A(net214),
    .X(instr_addr_o[23]));
 sky130_fd_sc_hd__buf_1 output210 (.A(net215),
    .X(instr_addr_o[24]));
 sky130_fd_sc_hd__buf_1 output211 (.A(net216),
    .X(instr_addr_o[25]));
 sky130_fd_sc_hd__buf_1 output212 (.A(net217),
    .X(instr_addr_o[26]));
 sky130_fd_sc_hd__buf_1 output213 (.A(net218),
    .X(instr_addr_o[27]));
 sky130_fd_sc_hd__buf_1 output214 (.A(net219),
    .X(instr_addr_o[28]));
 sky130_fd_sc_hd__buf_1 output215 (.A(net220),
    .X(instr_addr_o[29]));
 sky130_fd_sc_hd__buf_1 output216 (.A(net221),
    .X(instr_addr_o[2]));
 sky130_fd_sc_hd__buf_1 output217 (.A(net222),
    .X(instr_addr_o[30]));
 sky130_fd_sc_hd__buf_1 output218 (.A(net223),
    .X(instr_addr_o[31]));
 sky130_fd_sc_hd__buf_1 output219 (.A(net224),
    .X(instr_addr_o[3]));
 sky130_fd_sc_hd__buf_1 output220 (.A(net225),
    .X(instr_addr_o[4]));
 sky130_fd_sc_hd__buf_1 output221 (.A(net226),
    .X(instr_addr_o[5]));
 sky130_fd_sc_hd__buf_1 output222 (.A(net227),
    .X(instr_addr_o[6]));
 sky130_fd_sc_hd__buf_1 output223 (.A(net228),
    .X(instr_addr_o[7]));
 sky130_fd_sc_hd__buf_1 output224 (.A(net229),
    .X(instr_addr_o[8]));
 sky130_fd_sc_hd__buf_1 output225 (.A(net230),
    .X(instr_addr_o[9]));
 sky130_fd_sc_hd__buf_1 output226 (.A(net231),
    .X(instr_fetch_err_o));
 sky130_fd_sc_hd__buf_1 output227 (.A(net232),
    .X(instr_fetch_err_plus2_o));
 sky130_fd_sc_hd__buf_1 output228 (.A(net233),
    .X(instr_is_compressed_id_o));
 sky130_fd_sc_hd__buf_1 output229 (.A(net234),
    .X(instr_new_id_o));
 sky130_fd_sc_hd__buf_1 output230 (.A(net235),
    .X(instr_rdata_alu_id_o[0]));
 sky130_fd_sc_hd__buf_1 output231 (.A(net236),
    .X(instr_rdata_alu_id_o[10]));
 sky130_fd_sc_hd__buf_1 output232 (.A(net237),
    .X(instr_rdata_alu_id_o[11]));
 sky130_fd_sc_hd__buf_1 output233 (.A(net238),
    .X(instr_rdata_alu_id_o[12]));
 sky130_fd_sc_hd__buf_1 output234 (.A(net239),
    .X(instr_rdata_alu_id_o[13]));
 sky130_fd_sc_hd__buf_1 output235 (.A(net240),
    .X(instr_rdata_alu_id_o[14]));
 sky130_fd_sc_hd__buf_1 output236 (.A(net241),
    .X(instr_rdata_alu_id_o[15]));
 sky130_fd_sc_hd__buf_1 output237 (.A(net242),
    .X(instr_rdata_alu_id_o[16]));
 sky130_fd_sc_hd__buf_1 output238 (.A(net243),
    .X(instr_rdata_alu_id_o[17]));
 sky130_fd_sc_hd__buf_1 output239 (.A(net244),
    .X(instr_rdata_alu_id_o[18]));
 sky130_fd_sc_hd__buf_1 output240 (.A(net245),
    .X(instr_rdata_alu_id_o[19]));
 sky130_fd_sc_hd__buf_1 output241 (.A(net246),
    .X(instr_rdata_alu_id_o[1]));
 sky130_fd_sc_hd__buf_1 output242 (.A(net247),
    .X(instr_rdata_alu_id_o[20]));
 sky130_fd_sc_hd__buf_1 output243 (.A(net248),
    .X(instr_rdata_alu_id_o[21]));
 sky130_fd_sc_hd__buf_1 output244 (.A(net249),
    .X(instr_rdata_alu_id_o[22]));
 sky130_fd_sc_hd__buf_1 output245 (.A(net250),
    .X(instr_rdata_alu_id_o[23]));
 sky130_fd_sc_hd__buf_1 output246 (.A(net251),
    .X(instr_rdata_alu_id_o[24]));
 sky130_fd_sc_hd__buf_1 output247 (.A(net252),
    .X(instr_rdata_alu_id_o[25]));
 sky130_fd_sc_hd__buf_1 output248 (.A(net253),
    .X(instr_rdata_alu_id_o[26]));
 sky130_fd_sc_hd__buf_1 output249 (.A(net254),
    .X(instr_rdata_alu_id_o[27]));
 sky130_fd_sc_hd__buf_1 output250 (.A(net255),
    .X(instr_rdata_alu_id_o[28]));
 sky130_fd_sc_hd__buf_1 output251 (.A(net256),
    .X(instr_rdata_alu_id_o[29]));
 sky130_fd_sc_hd__buf_1 output252 (.A(net257),
    .X(instr_rdata_alu_id_o[2]));
 sky130_fd_sc_hd__buf_1 output253 (.A(net258),
    .X(instr_rdata_alu_id_o[30]));
 sky130_fd_sc_hd__buf_1 output254 (.A(net259),
    .X(instr_rdata_alu_id_o[31]));
 sky130_fd_sc_hd__buf_1 output255 (.A(net260),
    .X(instr_rdata_alu_id_o[3]));
 sky130_fd_sc_hd__buf_1 output256 (.A(net261),
    .X(instr_rdata_alu_id_o[4]));
 sky130_fd_sc_hd__buf_1 output257 (.A(net262),
    .X(instr_rdata_alu_id_o[5]));
 sky130_fd_sc_hd__buf_1 output258 (.A(net263),
    .X(instr_rdata_alu_id_o[6]));
 sky130_fd_sc_hd__buf_1 output259 (.A(net264),
    .X(instr_rdata_alu_id_o[7]));
 sky130_fd_sc_hd__buf_1 output260 (.A(net265),
    .X(instr_rdata_alu_id_o[8]));
 sky130_fd_sc_hd__buf_1 output261 (.A(net266),
    .X(instr_rdata_alu_id_o[9]));
 sky130_fd_sc_hd__buf_1 output262 (.A(net267),
    .X(instr_rdata_c_id_o[0]));
 sky130_fd_sc_hd__buf_1 output263 (.A(net268),
    .X(instr_rdata_c_id_o[10]));
 sky130_fd_sc_hd__buf_1 output264 (.A(net269),
    .X(instr_rdata_c_id_o[11]));
 sky130_fd_sc_hd__buf_1 output265 (.A(net270),
    .X(instr_rdata_c_id_o[12]));
 sky130_fd_sc_hd__buf_1 output266 (.A(net271),
    .X(instr_rdata_c_id_o[13]));
 sky130_fd_sc_hd__buf_1 output267 (.A(net272),
    .X(instr_rdata_c_id_o[14]));
 sky130_fd_sc_hd__buf_1 output268 (.A(net273),
    .X(instr_rdata_c_id_o[15]));
 sky130_fd_sc_hd__buf_1 output269 (.A(net274),
    .X(instr_rdata_c_id_o[1]));
 sky130_fd_sc_hd__buf_1 output270 (.A(net275),
    .X(instr_rdata_c_id_o[2]));
 sky130_fd_sc_hd__buf_1 output271 (.A(net276),
    .X(instr_rdata_c_id_o[3]));
 sky130_fd_sc_hd__buf_1 output272 (.A(net277),
    .X(instr_rdata_c_id_o[4]));
 sky130_fd_sc_hd__buf_1 output273 (.A(net278),
    .X(instr_rdata_c_id_o[5]));
 sky130_fd_sc_hd__buf_1 output274 (.A(net279),
    .X(instr_rdata_c_id_o[6]));
 sky130_fd_sc_hd__buf_1 output275 (.A(net280),
    .X(instr_rdata_c_id_o[7]));
 sky130_fd_sc_hd__buf_1 output276 (.A(net281),
    .X(instr_rdata_c_id_o[8]));
 sky130_fd_sc_hd__buf_1 output277 (.A(net282),
    .X(instr_rdata_c_id_o[9]));
 sky130_fd_sc_hd__buf_1 output278 (.A(net283),
    .X(instr_rdata_id_o[0]));
 sky130_fd_sc_hd__buf_1 output279 (.A(net284),
    .X(instr_rdata_id_o[10]));
 sky130_fd_sc_hd__buf_1 output280 (.A(net285),
    .X(instr_rdata_id_o[11]));
 sky130_fd_sc_hd__buf_1 output281 (.A(net286),
    .X(instr_rdata_id_o[12]));
 sky130_fd_sc_hd__buf_1 output282 (.A(net287),
    .X(instr_rdata_id_o[13]));
 sky130_fd_sc_hd__buf_1 output283 (.A(net288),
    .X(instr_rdata_id_o[14]));
 sky130_fd_sc_hd__buf_1 output284 (.A(net289),
    .X(instr_rdata_id_o[15]));
 sky130_fd_sc_hd__buf_1 output285 (.A(net290),
    .X(instr_rdata_id_o[16]));
 sky130_fd_sc_hd__buf_1 output286 (.A(net291),
    .X(instr_rdata_id_o[17]));
 sky130_fd_sc_hd__buf_1 output287 (.A(net292),
    .X(instr_rdata_id_o[18]));
 sky130_fd_sc_hd__buf_1 output288 (.A(net293),
    .X(instr_rdata_id_o[19]));
 sky130_fd_sc_hd__buf_1 output289 (.A(net294),
    .X(instr_rdata_id_o[1]));
 sky130_fd_sc_hd__buf_1 output290 (.A(net295),
    .X(instr_rdata_id_o[20]));
 sky130_fd_sc_hd__buf_1 output291 (.A(net296),
    .X(instr_rdata_id_o[21]));
 sky130_fd_sc_hd__buf_1 output292 (.A(net297),
    .X(instr_rdata_id_o[22]));
 sky130_fd_sc_hd__buf_1 output293 (.A(net298),
    .X(instr_rdata_id_o[23]));
 sky130_fd_sc_hd__buf_1 output294 (.A(net299),
    .X(instr_rdata_id_o[24]));
 sky130_fd_sc_hd__buf_1 output295 (.A(net300),
    .X(instr_rdata_id_o[25]));
 sky130_fd_sc_hd__buf_1 output296 (.A(net301),
    .X(instr_rdata_id_o[26]));
 sky130_fd_sc_hd__buf_1 output297 (.A(net302),
    .X(instr_rdata_id_o[27]));
 sky130_fd_sc_hd__buf_1 output298 (.A(net303),
    .X(instr_rdata_id_o[28]));
 sky130_fd_sc_hd__buf_1 output299 (.A(net304),
    .X(instr_rdata_id_o[29]));
 sky130_fd_sc_hd__buf_1 output300 (.A(net305),
    .X(instr_rdata_id_o[2]));
 sky130_fd_sc_hd__buf_1 output301 (.A(net306),
    .X(instr_rdata_id_o[30]));
 sky130_fd_sc_hd__buf_1 output302 (.A(net307),
    .X(instr_rdata_id_o[31]));
 sky130_fd_sc_hd__buf_1 output303 (.A(net308),
    .X(instr_rdata_id_o[3]));
 sky130_fd_sc_hd__buf_1 output304 (.A(net309),
    .X(instr_rdata_id_o[4]));
 sky130_fd_sc_hd__buf_1 output305 (.A(net310),
    .X(instr_rdata_id_o[5]));
 sky130_fd_sc_hd__buf_1 output306 (.A(net311),
    .X(instr_rdata_id_o[6]));
 sky130_fd_sc_hd__buf_1 output307 (.A(net312),
    .X(instr_rdata_id_o[7]));
 sky130_fd_sc_hd__buf_1 output308 (.A(net313),
    .X(instr_rdata_id_o[8]));
 sky130_fd_sc_hd__buf_1 output309 (.A(net314),
    .X(instr_rdata_id_o[9]));
 sky130_fd_sc_hd__buf_1 output310 (.A(net315),
    .X(instr_req_o));
 sky130_fd_sc_hd__buf_1 output311 (.A(net316),
    .X(instr_valid_id_o));
 sky130_fd_sc_hd__buf_1 output312 (.A(net317),
    .X(pc_id_o[10]));
 sky130_fd_sc_hd__buf_1 output313 (.A(net318),
    .X(pc_id_o[11]));
 sky130_fd_sc_hd__buf_1 output314 (.A(net319),
    .X(pc_id_o[12]));
 sky130_fd_sc_hd__buf_1 output315 (.A(net320),
    .X(pc_id_o[13]));
 sky130_fd_sc_hd__buf_1 output316 (.A(net321),
    .X(pc_id_o[14]));
 sky130_fd_sc_hd__buf_1 output317 (.A(net322),
    .X(pc_id_o[15]));
 sky130_fd_sc_hd__buf_1 output318 (.A(net323),
    .X(pc_id_o[16]));
 sky130_fd_sc_hd__buf_1 output319 (.A(net324),
    .X(pc_id_o[17]));
 sky130_fd_sc_hd__buf_1 output320 (.A(net325),
    .X(pc_id_o[18]));
 sky130_fd_sc_hd__buf_1 output321 (.A(net326),
    .X(pc_id_o[19]));
 sky130_fd_sc_hd__buf_1 output322 (.A(net327),
    .X(pc_id_o[1]));
 sky130_fd_sc_hd__buf_1 output323 (.A(net328),
    .X(pc_id_o[20]));
 sky130_fd_sc_hd__buf_1 output324 (.A(net329),
    .X(pc_id_o[21]));
 sky130_fd_sc_hd__buf_1 output325 (.A(net330),
    .X(pc_id_o[22]));
 sky130_fd_sc_hd__buf_1 output326 (.A(net331),
    .X(pc_id_o[23]));
 sky130_fd_sc_hd__buf_1 output327 (.A(net332),
    .X(pc_id_o[24]));
 sky130_fd_sc_hd__buf_1 output328 (.A(net333),
    .X(pc_id_o[25]));
 sky130_fd_sc_hd__buf_1 output329 (.A(net334),
    .X(pc_id_o[26]));
 sky130_fd_sc_hd__buf_1 output330 (.A(net335),
    .X(pc_id_o[27]));
 sky130_fd_sc_hd__buf_1 output331 (.A(net336),
    .X(pc_id_o[28]));
 sky130_fd_sc_hd__buf_1 output332 (.A(net337),
    .X(pc_id_o[29]));
 sky130_fd_sc_hd__buf_1 output333 (.A(net338),
    .X(pc_id_o[2]));
 sky130_fd_sc_hd__buf_1 output334 (.A(net339),
    .X(pc_id_o[30]));
 sky130_fd_sc_hd__buf_1 output335 (.A(net340),
    .X(pc_id_o[31]));
 sky130_fd_sc_hd__buf_1 output336 (.A(net341),
    .X(pc_id_o[3]));
 sky130_fd_sc_hd__buf_1 output337 (.A(net342),
    .X(pc_id_o[4]));
 sky130_fd_sc_hd__buf_1 output338 (.A(net343),
    .X(pc_id_o[5]));
 sky130_fd_sc_hd__buf_1 output339 (.A(net344),
    .X(pc_id_o[6]));
 sky130_fd_sc_hd__buf_1 output340 (.A(net345),
    .X(pc_id_o[7]));
 sky130_fd_sc_hd__buf_1 output341 (.A(net346),
    .X(pc_id_o[8]));
 sky130_fd_sc_hd__buf_1 output342 (.A(net347),
    .X(pc_id_o[9]));
 sky130_fd_sc_hd__buf_1 output343 (.A(net348),
    .X(pc_if_o[10]));
 sky130_fd_sc_hd__buf_1 output344 (.A(net349),
    .X(pc_if_o[11]));
 sky130_fd_sc_hd__buf_1 output345 (.A(net350),
    .X(pc_if_o[12]));
 sky130_fd_sc_hd__buf_1 output346 (.A(net351),
    .X(pc_if_o[13]));
 sky130_fd_sc_hd__buf_1 output347 (.A(net352),
    .X(pc_if_o[14]));
 sky130_fd_sc_hd__buf_1 output348 (.A(net353),
    .X(pc_if_o[15]));
 sky130_fd_sc_hd__buf_1 output349 (.A(net354),
    .X(pc_if_o[16]));
 sky130_fd_sc_hd__buf_1 output350 (.A(net355),
    .X(pc_if_o[17]));
 sky130_fd_sc_hd__buf_1 output351 (.A(net356),
    .X(pc_if_o[18]));
 sky130_fd_sc_hd__buf_1 output352 (.A(net357),
    .X(pc_if_o[19]));
 sky130_fd_sc_hd__buf_1 output353 (.A(net358),
    .X(pc_if_o[1]));
 sky130_fd_sc_hd__buf_1 output354 (.A(net359),
    .X(pc_if_o[20]));
 sky130_fd_sc_hd__buf_1 output355 (.A(net360),
    .X(pc_if_o[21]));
 sky130_fd_sc_hd__buf_1 output356 (.A(net361),
    .X(pc_if_o[22]));
 sky130_fd_sc_hd__buf_1 output357 (.A(net362),
    .X(pc_if_o[23]));
 sky130_fd_sc_hd__buf_1 output358 (.A(net363),
    .X(pc_if_o[24]));
 sky130_fd_sc_hd__buf_1 output359 (.A(net364),
    .X(pc_if_o[25]));
 sky130_fd_sc_hd__buf_1 output360 (.A(net365),
    .X(pc_if_o[26]));
 sky130_fd_sc_hd__buf_1 output361 (.A(net366),
    .X(pc_if_o[27]));
 sky130_fd_sc_hd__buf_1 output362 (.A(net367),
    .X(pc_if_o[28]));
 sky130_fd_sc_hd__buf_1 output363 (.A(net368),
    .X(pc_if_o[29]));
 sky130_fd_sc_hd__buf_1 output364 (.A(net369),
    .X(pc_if_o[2]));
 sky130_fd_sc_hd__buf_1 output365 (.A(net370),
    .X(pc_if_o[30]));
 sky130_fd_sc_hd__buf_1 output366 (.A(net371),
    .X(pc_if_o[31]));
 sky130_fd_sc_hd__buf_1 output367 (.A(net372),
    .X(pc_if_o[3]));
 sky130_fd_sc_hd__buf_1 output368 (.A(net373),
    .X(pc_if_o[4]));
 sky130_fd_sc_hd__buf_1 output369 (.A(net374),
    .X(pc_if_o[5]));
 sky130_fd_sc_hd__buf_1 output370 (.A(net375),
    .X(pc_if_o[6]));
 sky130_fd_sc_hd__buf_1 output371 (.A(net376),
    .X(pc_if_o[7]));
 sky130_fd_sc_hd__buf_1 output372 (.A(net377),
    .X(pc_if_o[8]));
 sky130_fd_sc_hd__buf_1 output373 (.A(net378),
    .X(pc_if_o[9]));
 sky130_fd_sc_hd__conb_1 _2366__374 (.LO(net379));
 sky130_fd_sc_hd__conb_1 _2367__375 (.LO(net380));
 sky130_fd_sc_hd__conb_1 _2368__376 (.LO(net381));
 sky130_fd_sc_hd__conb_1 _2369__377 (.LO(net382));
 sky130_fd_sc_hd__conb_1 _2402__378 (.LO(net383));
 sky130_fd_sc_hd__conb_1 _2403__379 (.LO(net384));
 sky130_fd_sc_hd__conb_1 _2404__380 (.LO(net385));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk_i (.A(clknet_2_0__leaf_clk_i),
    .X(clknet_leaf_1_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk_i (.A(clknet_2_0__leaf_clk_i),
    .X(clknet_leaf_2_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk_i (.A(clknet_2_0__leaf_clk_i),
    .X(clknet_leaf_3_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk_i (.A(clknet_2_1__leaf_clk_i),
    .X(clknet_leaf_4_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk_i (.A(clknet_2_1__leaf_clk_i),
    .X(clknet_leaf_5_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk_i (.A(clknet_2_1__leaf_clk_i),
    .X(clknet_leaf_6_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk_i (.A(clknet_2_1__leaf_clk_i),
    .X(clknet_leaf_7_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk_i (.A(clknet_2_1__leaf_clk_i),
    .X(clknet_leaf_8_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk_i (.A(clknet_2_1__leaf_clk_i),
    .X(clknet_leaf_9_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk_i (.A(clknet_2_3__leaf_clk_i),
    .X(clknet_leaf_10_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk_i (.A(clknet_2_3__leaf_clk_i),
    .X(clknet_leaf_11_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk_i (.A(clknet_2_3__leaf_clk_i),
    .X(clknet_leaf_12_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk_i (.A(clknet_2_3__leaf_clk_i),
    .X(clknet_leaf_13_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk_i (.A(clknet_2_3__leaf_clk_i),
    .X(clknet_leaf_14_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk_i (.A(clknet_2_3__leaf_clk_i),
    .X(clknet_leaf_15_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk_i (.A(clknet_2_3__leaf_clk_i),
    .X(clknet_leaf_16_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk_i (.A(clknet_2_3__leaf_clk_i),
    .X(clknet_leaf_17_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk_i (.A(clknet_2_2__leaf_clk_i),
    .X(clknet_leaf_18_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk_i (.A(clknet_2_2__leaf_clk_i),
    .X(clknet_leaf_19_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk_i (.A(clknet_2_2__leaf_clk_i),
    .X(clknet_leaf_20_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk_i (.A(clknet_2_2__leaf_clk_i),
    .X(clknet_leaf_21_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk_i (.A(clknet_2_2__leaf_clk_i),
    .X(clknet_leaf_22_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk_i (.A(clknet_2_2__leaf_clk_i),
    .X(clknet_leaf_23_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk_i (.A(clknet_2_2__leaf_clk_i),
    .X(clknet_leaf_24_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk_i (.A(clknet_2_2__leaf_clk_i),
    .X(clknet_leaf_25_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk_i (.A(clknet_2_2__leaf_clk_i),
    .X(clknet_leaf_26_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk_i (.A(clknet_2_2__leaf_clk_i),
    .X(clknet_leaf_27_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk_i (.A(clknet_2_2__leaf_clk_i),
    .X(clknet_leaf_28_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk_i (.A(clknet_2_2__leaf_clk_i),
    .X(clknet_leaf_29_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk_i (.A(clknet_2_0__leaf_clk_i),
    .X(clknet_leaf_30_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk_i (.A(clknet_2_2__leaf_clk_i),
    .X(clknet_leaf_31_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk_i (.A(clknet_2_0__leaf_clk_i),
    .X(clknet_leaf_32_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk_i (.A(clknet_2_0__leaf_clk_i),
    .X(clknet_leaf_33_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk_i (.A(clknet_2_0__leaf_clk_i),
    .X(clknet_leaf_34_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk_i (.A(clk_i),
    .X(clknet_0_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_2_0__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_2_1__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_2_2__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_2_3__leaf_clk_i));
 sky130_fd_sc_hd__clkinv_16 clkload0 (.A(clknet_2_0__leaf_clk_i));
 sky130_fd_sc_hd__clkinv_16 clkload1 (.A(clknet_2_1__leaf_clk_i));
 sky130_fd_sc_hd__clkinv_16 clkload2 (.A(clknet_2_3__leaf_clk_i));
 sky130_fd_sc_hd__clkinv_1 clkload3 (.A(clknet_leaf_0_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkload4 (.A(clknet_leaf_1_clk_i));
 sky130_fd_sc_hd__clkinv_2 clkload5 (.A(clknet_leaf_2_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkload6 (.A(clknet_leaf_3_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkload7 (.A(clknet_leaf_30_clk_i));
 sky130_fd_sc_hd__clkinv_1 clkload8 (.A(clknet_leaf_32_clk_i));
 sky130_fd_sc_hd__clkinv_4 clkload9 (.A(clknet_leaf_34_clk_i));
 sky130_fd_sc_hd__bufinv_16 clkload10 (.A(clknet_leaf_5_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkload11 (.A(clknet_leaf_6_clk_i));
 sky130_fd_sc_hd__clkinv_1 clkload12 (.A(clknet_leaf_7_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkload13 (.A(clknet_leaf_8_clk_i));
 sky130_fd_sc_hd__inv_6 clkload14 (.A(clknet_leaf_18_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkload15 (.A(clknet_leaf_19_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkload16 (.A(clknet_leaf_20_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkload17 (.A(clknet_leaf_21_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkload18 (.A(clknet_leaf_22_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkload19 (.A(clknet_leaf_23_clk_i));
 sky130_fd_sc_hd__clkinv_2 clkload20 (.A(clknet_leaf_24_clk_i));
 sky130_fd_sc_hd__clkbuf_1 clkload21 (.A(clknet_leaf_25_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkload22 (.A(clknet_leaf_26_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkload23 (.A(clknet_leaf_27_clk_i));
 sky130_fd_sc_hd__clkinv_2 clkload24 (.A(clknet_leaf_28_clk_i));
 sky130_fd_sc_hd__clkinv_1 clkload25 (.A(clknet_leaf_31_clk_i));
 sky130_fd_sc_hd__clkinv_1 clkload26 (.A(clknet_leaf_11_clk_i));
 sky130_fd_sc_hd__clkinvlp_4 clkload27 (.A(clknet_leaf_12_clk_i));
 sky130_fd_sc_hd__clkinvlp_4 clkload28 (.A(clknet_leaf_13_clk_i));
 sky130_fd_sc_hd__clkinv_1 clkload29 (.A(clknet_leaf_14_clk_i));
 sky130_fd_sc_hd__clkinv_2 clkload30 (.A(clknet_leaf_15_clk_i));
 sky130_fd_sc_hd__clkinvlp_4 clkload31 (.A(clknet_leaf_16_clk_i));
 sky130_fd_sc_hd__clkinvlp_4 clkload32 (.A(clknet_leaf_17_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(net3));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_356 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_438 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_469 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_473 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_487 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_252 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_260 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_276 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_383 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_411 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_529 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_625 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_487 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_495 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_535 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_586 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_594 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_602 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_610 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_618 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_626 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_507 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_555 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_567 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_625 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_478 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_560 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_625 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_442 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_520 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_528 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_544 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_560 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_516 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_524 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_560 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_576 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_625 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_355 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_591 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_325 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_396 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_567 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_625 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_423 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_431 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_543 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_555 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_336 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_455 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_518 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_574 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_536 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_325 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_397 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_624 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_636 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_283 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_294 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_396 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_502 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_514 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_612 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_620 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_636 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_475 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_531 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_547 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_555 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_487 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_522 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_528 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_619 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_366 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_380 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_453 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_568 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_586 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_594 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_602 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_610 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_618 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_626 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_387 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_438 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_463 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_517 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_564 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_572 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_580 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_588 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_616 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_319 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_494 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_618 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_626 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_273 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_308 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_319 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_438 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_454 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_516 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_524 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_522 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_530 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_270 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_306 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_319 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_327 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_370 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_378 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_394 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_402 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_453 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_516 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_524 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_576 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_621 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_375 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_425 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_486 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_494 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_502 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_517 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_535 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_547 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_580 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_588 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_596 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_610 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_622 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_378 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_394 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_410 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_453 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_560 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_625 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_290 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_306 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_454 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_462 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_435 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_590 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_106 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_114 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_122 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_187 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_234 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_252 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_302 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_306 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_366 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_380 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_550 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_622 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_79 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_363 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_406 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_550 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_558 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_574 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_627 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_200 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_242 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_286 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_294 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_302 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_326 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_397 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_548 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_556 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_83 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_90 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_171 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_183 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_200 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_319 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_442 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_499 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_507 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_546 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_550 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_311 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_319 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_402 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_410 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_438 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_600 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_276 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_443 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_625 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_634 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_184 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_415 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_470 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_486 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_494 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_292 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_305 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_12 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_190 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_402 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_547 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_325 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_441 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_456 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_512 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_520 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_528 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_536 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_576 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_357 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_438 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_595 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_610 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_618 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_514 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_522 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_565 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_625 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_142 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_186 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_244 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_252 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_273 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_487 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_495 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_530 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_546 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_562 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_83 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_139 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_147 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_517 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_528 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_536 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_6 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_20 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_86 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_122 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_206 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_217 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_228 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_244 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_252 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_427 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_469 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_492 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_500 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_562 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_75 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_83 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_140 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_375 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_392 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_478 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_535 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_558 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_563 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_625 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_206 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_228 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_244 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_252 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_363 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_375 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_414 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_468 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_606 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_75 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_79 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_87 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_156 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_375 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_472 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_517 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_558 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_574 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_624 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_7 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_426 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_434 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_442 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_466 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_474 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_482 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_490 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_498 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_542 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_555 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_212 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_441 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_522 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_531 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_620 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_636 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_79 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_252 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_427 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_531 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_634 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_7 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_141 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_203 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_267 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_435 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_518 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_530 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_558 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_574 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_621 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_630 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_187 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_199 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_306 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_410 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_426 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_471 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_486 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_495 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_7 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_38 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_270 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_425 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_507 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_556 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_563 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_217 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_237 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_306 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_430 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_471 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_487 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_6 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_50 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_494 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_507 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_559 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_567 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_625 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_51 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_70 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_140 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_228 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_244 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_295 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_415 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_204 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_342 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_390 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_406 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_432 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_469 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_514 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_522 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_534 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_576 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_592 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_273 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_283 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_319 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_413 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_462 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_470 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_486 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_502 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_524 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_530 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_546 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_52 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_203 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_321 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_396 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_456 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_503 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_512 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_520 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_536 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_563 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_619 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_60 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_186 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_295 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_415 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_427 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_469 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_495 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_562 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_618 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_626 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_40 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_290 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_315 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_323 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_550 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_558 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_574 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_624 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_74 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_295 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_490 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_498 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_535 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_78 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_112 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_207 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_267 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_441 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_454 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_503 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_514 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_525 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_411 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_453 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_460 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_522 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_530 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_595 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_607 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_76 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_84 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_92 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_154 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_248 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_342 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_392 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_404 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_528 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_624 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_201 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_234 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_411 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_441 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_530 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_561 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_90 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_193 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_210 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_483 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_506 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_7 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_15 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_422 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_524 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_530 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_546 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_622 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_13 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_340 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_438 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_446 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_529 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_560 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_621 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_214 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_222 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_236 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_244 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_405 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_420 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_428 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_448 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_472 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_480 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_487 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_495 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_526 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_534 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_542 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_623 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_223 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_231 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_276 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_413 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_453 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_488 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_517 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_627 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_634 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_6 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_170 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_186 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_291 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_364 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_372 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_415 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_528 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_544 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_595 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_612 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_234 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_264 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_452 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_462 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_478 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_503 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_516 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_562 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_570 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_578 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_586 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_246 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_415 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_502 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_524 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_530 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_595 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_610 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_618 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_94 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_210 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_427 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_470 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_501 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_522 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_605 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_46 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_54 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_70 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_78 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_306 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_366 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_374 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_428 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_468 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_484 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_492 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_504 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_522 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_540 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_548 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_560 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_612 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_191 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_264 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_303 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_315 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_323 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_453 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_517 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_630 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_33 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_182 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_206 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_528 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_544 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_603 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_637 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_20 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_140 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_207 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_330 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_439 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_447 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_495 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_564 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_572 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_580 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_588 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_618 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_634 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_46 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_54 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_62 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_113 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_156 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_180 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_247 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_291 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_357 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_439 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_466 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_471 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_487 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_495 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_516 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_531 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_634 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_80 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_393 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_440 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_512 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_524 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_575 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_605 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_630 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_111 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_246 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_351 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_375 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_428 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_515 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_11 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_23 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_54 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_160 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_216 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_251 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_276 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_292 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_575 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_610 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_618 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_634 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_192 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_446 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_480 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_488 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_40 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_193 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_321 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_441 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_585 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_616 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_624 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_375 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_425 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_492 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_590 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_602 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_637 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_70 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_83 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_454 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_468 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_567 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_625 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_183 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_424 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_432 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_498 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_562 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_590 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_606 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_21 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_166 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_202 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_222 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_252 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_260 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_312 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_324 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_342 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_622 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_127 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_139 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_201 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_274 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_302 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_323 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_366 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_374 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_491 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_531 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_556 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_90 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_98 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_402 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_514 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_574 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_625 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_637 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_174 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_182 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_357 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_550 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_595 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_619 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_634 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_70 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_79 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_87 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_103 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_210 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_236 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_246 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_375 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_625 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_595 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_605 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_618 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_626 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_634 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_180 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_226 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_231 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_84 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_150 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_207 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_228 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_232 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_251 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_321 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_625 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_7 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_15 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_70 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_123 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_595 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_618 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_626 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_637 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_25 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_66 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_92 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_191 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_251 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_303 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_610 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_618 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_626 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_634 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_70 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_180 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_337 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_362 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_595 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_196 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_204 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_212 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_623 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_108 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_186 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_5 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_13 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_21 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_152 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_212 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_610 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_618 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_626 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_634 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_170 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_182 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_357 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_595 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_5 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_13 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_21 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_220 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_625 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_321 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_463 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_471 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_487 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_495 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_603 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_435 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_440 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_456 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_500 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_522 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_581 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_626 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_634 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_10 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_20 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_86 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_170 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_247 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_259 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_303 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_565 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_623 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_637 ();
endmodule
