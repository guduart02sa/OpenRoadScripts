VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 1000 ;
END UNITS

VIA ibex_id_stage_via2_3_1600_480_1_5_320_320
  VIARULE M1M2_PR ;
  CUTSIZE 0.15 0.15 ;
  LAYERS met1 via met2 ;
  CUTSPACING 0.17 0.17 ;
  ENCLOSURE 0.085 0.165 0.055 0.085 ;
  ROWCOL 1 5 ;
END ibex_id_stage_via2_3_1600_480_1_5_320_320

VIA ibex_id_stage_via3_4_1600_480_1_4_400_400
  VIARULE M2M3_PR ;
  CUTSIZE 0.2 0.2 ;
  LAYERS met2 via2 met3 ;
  CUTSPACING 0.2 0.2 ;
  ENCLOSURE 0.04 0.085 0.065 0.065 ;
  ROWCOL 1 4 ;
END ibex_id_stage_via3_4_1600_480_1_4_400_400

VIA ibex_id_stage_via4_5_1600_480_1_4_400_400
  VIARULE M3M4_PR ;
  CUTSIZE 0.2 0.2 ;
  LAYERS met3 via3 met4 ;
  CUTSPACING 0.2 0.2 ;
  ENCLOSURE 0.09 0.06 0.1 0.065 ;
  ROWCOL 1 4 ;
END ibex_id_stage_via4_5_1600_480_1_4_400_400

VIA ibex_id_stage_via5_6_1600_1600_1_1_1600_1600
  VIARULE M4M5_PR ;
  CUTSIZE 0.8 0.8 ;
  LAYERS met4 via4 met5 ;
  CUTSPACING 0.8 0.8 ;
  ENCLOSURE 0.4 0.19 0.31 0.4 ;
END ibex_id_stage_via5_6_1600_1600_1_1_1600_1600

MACRO ibex_id_stage
  FOREIGN ibex_id_stage 0 0 ;
  CLASS BLOCK ;
  SIZE 177.52 BY 704.07 ;
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      LAYER met5 ;
        RECT  27.72 681.92 165.02 683.52 ;
        RECT  27.72 654.72 165.02 656.32 ;
        RECT  27.72 627.52 165.02 629.12 ;
        RECT  27.72 600.32 165.02 601.92 ;
        RECT  27.72 573.12 165.02 574.72 ;
        RECT  27.72 545.92 165.02 547.52 ;
        RECT  27.72 518.72 165.02 520.32 ;
        RECT  27.72 491.52 165.02 493.12 ;
        RECT  27.72 464.32 165.02 465.92 ;
        RECT  27.72 437.12 165.02 438.72 ;
        RECT  27.72 409.92 165.02 411.52 ;
        RECT  27.72 382.72 165.02 384.32 ;
        RECT  27.72 355.52 165.02 357.12 ;
        RECT  27.72 328.32 165.02 329.92 ;
        RECT  27.72 301.12 165.02 302.72 ;
        RECT  27.72 273.92 165.02 275.52 ;
        RECT  27.72 246.72 165.02 248.32 ;
        RECT  27.72 219.52 165.02 221.12 ;
        RECT  27.72 192.32 165.02 193.92 ;
        RECT  27.72 165.12 165.02 166.72 ;
        RECT  27.72 137.92 165.02 139.52 ;
        RECT  27.72 110.72 165.02 112.32 ;
        RECT  27.72 83.52 165.02 85.12 ;
        RECT  27.72 56.32 165.02 57.92 ;
        RECT  27.72 29.12 165.02 30.72 ;
      LAYER met4 ;
        RECT  163.42 5.2 165.02 702 ;
        RECT  136.28 5.2 137.88 702 ;
        RECT  109.14 5.2 110.74 702 ;
        RECT  82 5.2 83.6 702 ;
        RECT  54.86 5.2 56.46 702 ;
        RECT  27.72 5.2 29.32 702 ;
      LAYER met1 ;
        RECT  1.38 701.52 176.18 702 ;
        RECT  1.38 696.08 176.18 696.56 ;
        RECT  1.38 690.64 176.18 691.12 ;
        RECT  1.38 685.2 176.18 685.68 ;
        RECT  1.38 679.76 176.18 680.24 ;
        RECT  1.38 674.32 176.18 674.8 ;
        RECT  1.38 668.88 176.18 669.36 ;
        RECT  1.38 663.44 176.18 663.92 ;
        RECT  1.38 658 176.18 658.48 ;
        RECT  1.38 652.56 176.18 653.04 ;
        RECT  1.38 647.12 176.18 647.6 ;
        RECT  1.38 641.68 176.18 642.16 ;
        RECT  1.38 636.24 176.18 636.72 ;
        RECT  1.38 630.8 176.18 631.28 ;
        RECT  1.38 625.36 176.18 625.84 ;
        RECT  1.38 619.92 176.18 620.4 ;
        RECT  1.38 614.48 176.18 614.96 ;
        RECT  1.38 609.04 176.18 609.52 ;
        RECT  1.38 603.6 176.18 604.08 ;
        RECT  1.38 598.16 176.18 598.64 ;
        RECT  1.38 592.72 176.18 593.2 ;
        RECT  1.38 587.28 176.18 587.76 ;
        RECT  1.38 581.84 176.18 582.32 ;
        RECT  1.38 576.4 176.18 576.88 ;
        RECT  1.38 570.96 176.18 571.44 ;
        RECT  1.38 565.52 176.18 566 ;
        RECT  1.38 560.08 176.18 560.56 ;
        RECT  1.38 554.64 176.18 555.12 ;
        RECT  1.38 549.2 176.18 549.68 ;
        RECT  1.38 543.76 176.18 544.24 ;
        RECT  1.38 538.32 176.18 538.8 ;
        RECT  1.38 532.88 176.18 533.36 ;
        RECT  1.38 527.44 176.18 527.92 ;
        RECT  1.38 522 176.18 522.48 ;
        RECT  1.38 516.56 176.18 517.04 ;
        RECT  1.38 511.12 176.18 511.6 ;
        RECT  1.38 505.68 176.18 506.16 ;
        RECT  1.38 500.24 176.18 500.72 ;
        RECT  1.38 494.8 176.18 495.28 ;
        RECT  1.38 489.36 176.18 489.84 ;
        RECT  1.38 483.92 176.18 484.4 ;
        RECT  1.38 478.48 176.18 478.96 ;
        RECT  1.38 473.04 176.18 473.52 ;
        RECT  1.38 467.6 176.18 468.08 ;
        RECT  1.38 462.16 176.18 462.64 ;
        RECT  1.38 456.72 176.18 457.2 ;
        RECT  1.38 451.28 176.18 451.76 ;
        RECT  1.38 445.84 176.18 446.32 ;
        RECT  1.38 440.4 176.18 440.88 ;
        RECT  1.38 434.96 176.18 435.44 ;
        RECT  1.38 429.52 176.18 430 ;
        RECT  1.38 424.08 176.18 424.56 ;
        RECT  1.38 418.64 176.18 419.12 ;
        RECT  1.38 413.2 176.18 413.68 ;
        RECT  1.38 407.76 176.18 408.24 ;
        RECT  1.38 402.32 176.18 402.8 ;
        RECT  1.38 396.88 176.18 397.36 ;
        RECT  1.38 391.44 176.18 391.92 ;
        RECT  1.38 386 176.18 386.48 ;
        RECT  1.38 380.56 176.18 381.04 ;
        RECT  1.38 375.12 176.18 375.6 ;
        RECT  1.38 369.68 176.18 370.16 ;
        RECT  1.38 364.24 176.18 364.72 ;
        RECT  1.38 358.8 176.18 359.28 ;
        RECT  1.38 353.36 176.18 353.84 ;
        RECT  1.38 347.92 176.18 348.4 ;
        RECT  1.38 342.48 176.18 342.96 ;
        RECT  1.38 337.04 176.18 337.52 ;
        RECT  1.38 331.6 176.18 332.08 ;
        RECT  1.38 326.16 176.18 326.64 ;
        RECT  1.38 320.72 176.18 321.2 ;
        RECT  1.38 315.28 176.18 315.76 ;
        RECT  1.38 309.84 176.18 310.32 ;
        RECT  1.38 304.4 176.18 304.88 ;
        RECT  1.38 298.96 176.18 299.44 ;
        RECT  1.38 293.52 176.18 294 ;
        RECT  1.38 288.08 176.18 288.56 ;
        RECT  1.38 282.64 176.18 283.12 ;
        RECT  1.38 277.2 176.18 277.68 ;
        RECT  1.38 271.76 176.18 272.24 ;
        RECT  1.38 266.32 176.18 266.8 ;
        RECT  1.38 260.88 176.18 261.36 ;
        RECT  1.38 255.44 176.18 255.92 ;
        RECT  1.38 250 176.18 250.48 ;
        RECT  1.38 244.56 176.18 245.04 ;
        RECT  1.38 239.12 176.18 239.6 ;
        RECT  1.38 233.68 176.18 234.16 ;
        RECT  1.38 228.24 176.18 228.72 ;
        RECT  1.38 222.8 176.18 223.28 ;
        RECT  1.38 217.36 176.18 217.84 ;
        RECT  1.38 211.92 176.18 212.4 ;
        RECT  1.38 206.48 176.18 206.96 ;
        RECT  1.38 201.04 176.18 201.52 ;
        RECT  1.38 195.6 176.18 196.08 ;
        RECT  1.38 190.16 176.18 190.64 ;
        RECT  1.38 184.72 176.18 185.2 ;
        RECT  1.38 179.28 176.18 179.76 ;
        RECT  1.38 173.84 176.18 174.32 ;
        RECT  1.38 168.4 176.18 168.88 ;
        RECT  1.38 162.96 176.18 163.44 ;
        RECT  1.38 157.52 176.18 158 ;
        RECT  1.38 152.08 176.18 152.56 ;
        RECT  1.38 146.64 176.18 147.12 ;
        RECT  1.38 141.2 176.18 141.68 ;
        RECT  1.38 135.76 176.18 136.24 ;
        RECT  1.38 130.32 176.18 130.8 ;
        RECT  1.38 124.88 176.18 125.36 ;
        RECT  1.38 119.44 176.18 119.92 ;
        RECT  1.38 114 176.18 114.48 ;
        RECT  1.38 108.56 176.18 109.04 ;
        RECT  1.38 103.12 176.18 103.6 ;
        RECT  1.38 97.68 176.18 98.16 ;
        RECT  1.38 92.24 176.18 92.72 ;
        RECT  1.38 86.8 176.18 87.28 ;
        RECT  1.38 81.36 176.18 81.84 ;
        RECT  1.38 75.92 176.18 76.4 ;
        RECT  1.38 70.48 176.18 70.96 ;
        RECT  1.38 65.04 176.18 65.52 ;
        RECT  1.38 59.6 176.18 60.08 ;
        RECT  1.38 54.16 176.18 54.64 ;
        RECT  1.38 48.72 176.18 49.2 ;
        RECT  1.38 43.28 176.18 43.76 ;
        RECT  1.38 37.84 176.18 38.32 ;
        RECT  1.38 32.4 176.18 32.88 ;
        RECT  1.38 26.96 176.18 27.44 ;
        RECT  1.38 21.52 176.18 22 ;
        RECT  1.38 16.08 176.18 16.56 ;
        RECT  1.38 10.64 176.18 11.12 ;
        RECT  1.38 5.2 176.18 5.68 ;
      VIA 164.22 682.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 655.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 628.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 601.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 573.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 546.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 519.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 492.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 465.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 437.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 410.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 383.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 356.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 329.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 301.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 274.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 247.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 220.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 193.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 165.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 138.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 111.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 84.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 57.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 164.22 29.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 682.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 655.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 628.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 601.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 573.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 546.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 519.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 492.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 465.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 437.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 410.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 383.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 356.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 329.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 301.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 274.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 247.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 220.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 193.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 165.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 138.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 111.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 84.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 57.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 137.08 29.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 682.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 655.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 628.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 601.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 573.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 546.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 519.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 492.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 465.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 437.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 410.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 383.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 356.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 329.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 301.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 274.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 247.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 220.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 193.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 165.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 138.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 111.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 84.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 57.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 109.94 29.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 682.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 655.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 628.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 601.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 573.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 546.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 519.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 492.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 465.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 437.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 410.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 383.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 356.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 329.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 301.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 274.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 247.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 220.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 193.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 165.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 138.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 111.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 84.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 57.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 82.8 29.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 682.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 655.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 628.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 601.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 573.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 546.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 519.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 492.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 465.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 437.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 410.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 383.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 356.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 329.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 301.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 274.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 247.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 220.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 193.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 165.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 138.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 111.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 84.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 57.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 55.66 29.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 682.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 655.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 628.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 601.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 573.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 546.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 519.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 492.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 465.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 437.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 410.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 383.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 356.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 329.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 301.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 274.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 247.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 220.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 193.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 165.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 138.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 111.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 84.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 57.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 28.52 29.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      LAYER met3 ;
        RECT  163.43 701.595 165.01 701.925 ;
      VIA 164.22 701.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 701.575 164.99 701.945 ;
      VIA 164.22 701.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 701.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 696.155 165.01 696.485 ;
      VIA 164.22 696.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 696.135 164.99 696.505 ;
      VIA 164.22 696.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 696.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 690.715 165.01 691.045 ;
      VIA 164.22 690.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 690.695 164.99 691.065 ;
      VIA 164.22 690.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 690.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 685.275 165.01 685.605 ;
      VIA 164.22 685.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 685.255 164.99 685.625 ;
      VIA 164.22 685.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 685.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 679.835 165.01 680.165 ;
      VIA 164.22 680 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 679.815 164.99 680.185 ;
      VIA 164.22 680 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 680 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 674.395 165.01 674.725 ;
      VIA 164.22 674.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 674.375 164.99 674.745 ;
      VIA 164.22 674.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 674.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 668.955 165.01 669.285 ;
      VIA 164.22 669.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 668.935 164.99 669.305 ;
      VIA 164.22 669.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 669.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 663.515 165.01 663.845 ;
      VIA 164.22 663.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 663.495 164.99 663.865 ;
      VIA 164.22 663.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 663.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 658.075 165.01 658.405 ;
      VIA 164.22 658.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 658.055 164.99 658.425 ;
      VIA 164.22 658.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 658.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 652.635 165.01 652.965 ;
      VIA 164.22 652.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 652.615 164.99 652.985 ;
      VIA 164.22 652.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 652.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 647.195 165.01 647.525 ;
      VIA 164.22 647.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 647.175 164.99 647.545 ;
      VIA 164.22 647.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 647.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 641.755 165.01 642.085 ;
      VIA 164.22 641.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 641.735 164.99 642.105 ;
      VIA 164.22 641.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 641.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 636.315 165.01 636.645 ;
      VIA 164.22 636.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 636.295 164.99 636.665 ;
      VIA 164.22 636.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 636.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 630.875 165.01 631.205 ;
      VIA 164.22 631.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 630.855 164.99 631.225 ;
      VIA 164.22 631.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 631.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 625.435 165.01 625.765 ;
      VIA 164.22 625.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 625.415 164.99 625.785 ;
      VIA 164.22 625.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 625.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 619.995 165.01 620.325 ;
      VIA 164.22 620.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 619.975 164.99 620.345 ;
      VIA 164.22 620.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 620.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 614.555 165.01 614.885 ;
      VIA 164.22 614.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 614.535 164.99 614.905 ;
      VIA 164.22 614.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 614.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 609.115 165.01 609.445 ;
      VIA 164.22 609.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 609.095 164.99 609.465 ;
      VIA 164.22 609.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 609.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 603.675 165.01 604.005 ;
      VIA 164.22 603.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 603.655 164.99 604.025 ;
      VIA 164.22 603.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 603.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 598.235 165.01 598.565 ;
      VIA 164.22 598.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 598.215 164.99 598.585 ;
      VIA 164.22 598.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 598.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 592.795 165.01 593.125 ;
      VIA 164.22 592.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 592.775 164.99 593.145 ;
      VIA 164.22 592.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 592.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 587.355 165.01 587.685 ;
      VIA 164.22 587.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 587.335 164.99 587.705 ;
      VIA 164.22 587.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 587.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 581.915 165.01 582.245 ;
      VIA 164.22 582.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 581.895 164.99 582.265 ;
      VIA 164.22 582.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 582.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 576.475 165.01 576.805 ;
      VIA 164.22 576.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 576.455 164.99 576.825 ;
      VIA 164.22 576.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 576.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 571.035 165.01 571.365 ;
      VIA 164.22 571.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 571.015 164.99 571.385 ;
      VIA 164.22 571.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 571.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 565.595 165.01 565.925 ;
      VIA 164.22 565.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 565.575 164.99 565.945 ;
      VIA 164.22 565.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 565.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 560.155 165.01 560.485 ;
      VIA 164.22 560.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 560.135 164.99 560.505 ;
      VIA 164.22 560.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 560.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 554.715 165.01 555.045 ;
      VIA 164.22 554.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 554.695 164.99 555.065 ;
      VIA 164.22 554.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 554.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 549.275 165.01 549.605 ;
      VIA 164.22 549.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 549.255 164.99 549.625 ;
      VIA 164.22 549.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 549.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 543.835 165.01 544.165 ;
      VIA 164.22 544 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 543.815 164.99 544.185 ;
      VIA 164.22 544 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 544 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 538.395 165.01 538.725 ;
      VIA 164.22 538.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 538.375 164.99 538.745 ;
      VIA 164.22 538.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 538.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 532.955 165.01 533.285 ;
      VIA 164.22 533.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 532.935 164.99 533.305 ;
      VIA 164.22 533.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 533.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 527.515 165.01 527.845 ;
      VIA 164.22 527.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 527.495 164.99 527.865 ;
      VIA 164.22 527.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 527.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 522.075 165.01 522.405 ;
      VIA 164.22 522.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 522.055 164.99 522.425 ;
      VIA 164.22 522.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 522.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 516.635 165.01 516.965 ;
      VIA 164.22 516.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 516.615 164.99 516.985 ;
      VIA 164.22 516.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 516.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 511.195 165.01 511.525 ;
      VIA 164.22 511.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 511.175 164.99 511.545 ;
      VIA 164.22 511.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 511.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 505.755 165.01 506.085 ;
      VIA 164.22 505.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 505.735 164.99 506.105 ;
      VIA 164.22 505.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 505.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 500.315 165.01 500.645 ;
      VIA 164.22 500.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 500.295 164.99 500.665 ;
      VIA 164.22 500.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 500.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 494.875 165.01 495.205 ;
      VIA 164.22 495.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 494.855 164.99 495.225 ;
      VIA 164.22 495.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 495.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 489.435 165.01 489.765 ;
      VIA 164.22 489.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 489.415 164.99 489.785 ;
      VIA 164.22 489.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 489.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 483.995 165.01 484.325 ;
      VIA 164.22 484.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 483.975 164.99 484.345 ;
      VIA 164.22 484.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 484.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 478.555 165.01 478.885 ;
      VIA 164.22 478.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 478.535 164.99 478.905 ;
      VIA 164.22 478.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 478.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 473.115 165.01 473.445 ;
      VIA 164.22 473.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 473.095 164.99 473.465 ;
      VIA 164.22 473.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 473.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 467.675 165.01 468.005 ;
      VIA 164.22 467.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 467.655 164.99 468.025 ;
      VIA 164.22 467.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 467.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 462.235 165.01 462.565 ;
      VIA 164.22 462.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 462.215 164.99 462.585 ;
      VIA 164.22 462.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 462.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 456.795 165.01 457.125 ;
      VIA 164.22 456.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 456.775 164.99 457.145 ;
      VIA 164.22 456.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 456.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 451.355 165.01 451.685 ;
      VIA 164.22 451.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 451.335 164.99 451.705 ;
      VIA 164.22 451.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 451.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 445.915 165.01 446.245 ;
      VIA 164.22 446.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 445.895 164.99 446.265 ;
      VIA 164.22 446.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 446.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 440.475 165.01 440.805 ;
      VIA 164.22 440.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 440.455 164.99 440.825 ;
      VIA 164.22 440.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 440.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 435.035 165.01 435.365 ;
      VIA 164.22 435.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 435.015 164.99 435.385 ;
      VIA 164.22 435.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 435.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 429.595 165.01 429.925 ;
      VIA 164.22 429.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 429.575 164.99 429.945 ;
      VIA 164.22 429.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 429.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 424.155 165.01 424.485 ;
      VIA 164.22 424.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 424.135 164.99 424.505 ;
      VIA 164.22 424.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 424.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 418.715 165.01 419.045 ;
      VIA 164.22 418.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 418.695 164.99 419.065 ;
      VIA 164.22 418.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 418.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 413.275 165.01 413.605 ;
      VIA 164.22 413.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 413.255 164.99 413.625 ;
      VIA 164.22 413.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 413.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 407.835 165.01 408.165 ;
      VIA 164.22 408 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 407.815 164.99 408.185 ;
      VIA 164.22 408 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 408 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 402.395 165.01 402.725 ;
      VIA 164.22 402.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 402.375 164.99 402.745 ;
      VIA 164.22 402.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 402.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 396.955 165.01 397.285 ;
      VIA 164.22 397.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 396.935 164.99 397.305 ;
      VIA 164.22 397.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 397.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 391.515 165.01 391.845 ;
      VIA 164.22 391.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 391.495 164.99 391.865 ;
      VIA 164.22 391.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 391.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 386.075 165.01 386.405 ;
      VIA 164.22 386.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 386.055 164.99 386.425 ;
      VIA 164.22 386.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 386.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 380.635 165.01 380.965 ;
      VIA 164.22 380.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 380.615 164.99 380.985 ;
      VIA 164.22 380.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 380.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 375.195 165.01 375.525 ;
      VIA 164.22 375.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 375.175 164.99 375.545 ;
      VIA 164.22 375.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 375.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 369.755 165.01 370.085 ;
      VIA 164.22 369.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 369.735 164.99 370.105 ;
      VIA 164.22 369.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 369.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 364.315 165.01 364.645 ;
      VIA 164.22 364.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 364.295 164.99 364.665 ;
      VIA 164.22 364.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 364.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 358.875 165.01 359.205 ;
      VIA 164.22 359.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 358.855 164.99 359.225 ;
      VIA 164.22 359.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 359.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 353.435 165.01 353.765 ;
      VIA 164.22 353.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 353.415 164.99 353.785 ;
      VIA 164.22 353.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 353.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 347.995 165.01 348.325 ;
      VIA 164.22 348.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 347.975 164.99 348.345 ;
      VIA 164.22 348.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 348.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 342.555 165.01 342.885 ;
      VIA 164.22 342.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 342.535 164.99 342.905 ;
      VIA 164.22 342.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 342.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 337.115 165.01 337.445 ;
      VIA 164.22 337.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 337.095 164.99 337.465 ;
      VIA 164.22 337.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 337.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 331.675 165.01 332.005 ;
      VIA 164.22 331.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 331.655 164.99 332.025 ;
      VIA 164.22 331.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 331.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 326.235 165.01 326.565 ;
      VIA 164.22 326.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 326.215 164.99 326.585 ;
      VIA 164.22 326.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 326.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 320.795 165.01 321.125 ;
      VIA 164.22 320.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 320.775 164.99 321.145 ;
      VIA 164.22 320.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 320.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 315.355 165.01 315.685 ;
      VIA 164.22 315.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 315.335 164.99 315.705 ;
      VIA 164.22 315.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 315.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 309.915 165.01 310.245 ;
      VIA 164.22 310.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 309.895 164.99 310.265 ;
      VIA 164.22 310.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 310.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 304.475 165.01 304.805 ;
      VIA 164.22 304.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 304.455 164.99 304.825 ;
      VIA 164.22 304.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 304.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 299.035 165.01 299.365 ;
      VIA 164.22 299.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 299.015 164.99 299.385 ;
      VIA 164.22 299.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 299.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 293.595 165.01 293.925 ;
      VIA 164.22 293.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 293.575 164.99 293.945 ;
      VIA 164.22 293.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 293.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 288.155 165.01 288.485 ;
      VIA 164.22 288.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 288.135 164.99 288.505 ;
      VIA 164.22 288.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 288.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 282.715 165.01 283.045 ;
      VIA 164.22 282.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 282.695 164.99 283.065 ;
      VIA 164.22 282.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 282.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 277.275 165.01 277.605 ;
      VIA 164.22 277.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 277.255 164.99 277.625 ;
      VIA 164.22 277.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 277.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 271.835 165.01 272.165 ;
      VIA 164.22 272 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 271.815 164.99 272.185 ;
      VIA 164.22 272 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 272 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 266.395 165.01 266.725 ;
      VIA 164.22 266.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 266.375 164.99 266.745 ;
      VIA 164.22 266.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 266.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 260.955 165.01 261.285 ;
      VIA 164.22 261.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 260.935 164.99 261.305 ;
      VIA 164.22 261.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 261.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 255.515 165.01 255.845 ;
      VIA 164.22 255.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 255.495 164.99 255.865 ;
      VIA 164.22 255.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 255.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 250.075 165.01 250.405 ;
      VIA 164.22 250.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 250.055 164.99 250.425 ;
      VIA 164.22 250.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 250.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 244.635 165.01 244.965 ;
      VIA 164.22 244.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 244.615 164.99 244.985 ;
      VIA 164.22 244.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 244.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 239.195 165.01 239.525 ;
      VIA 164.22 239.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 239.175 164.99 239.545 ;
      VIA 164.22 239.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 239.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 233.755 165.01 234.085 ;
      VIA 164.22 233.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 233.735 164.99 234.105 ;
      VIA 164.22 233.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 233.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 228.315 165.01 228.645 ;
      VIA 164.22 228.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 228.295 164.99 228.665 ;
      VIA 164.22 228.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 228.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 222.875 165.01 223.205 ;
      VIA 164.22 223.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 222.855 164.99 223.225 ;
      VIA 164.22 223.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 223.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 217.435 165.01 217.765 ;
      VIA 164.22 217.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 217.415 164.99 217.785 ;
      VIA 164.22 217.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 217.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 211.995 165.01 212.325 ;
      VIA 164.22 212.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 211.975 164.99 212.345 ;
      VIA 164.22 212.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 212.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 206.555 165.01 206.885 ;
      VIA 164.22 206.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 206.535 164.99 206.905 ;
      VIA 164.22 206.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 206.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 201.115 165.01 201.445 ;
      VIA 164.22 201.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 201.095 164.99 201.465 ;
      VIA 164.22 201.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 201.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 195.675 165.01 196.005 ;
      VIA 164.22 195.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 195.655 164.99 196.025 ;
      VIA 164.22 195.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 195.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 190.235 165.01 190.565 ;
      VIA 164.22 190.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 190.215 164.99 190.585 ;
      VIA 164.22 190.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 190.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 184.795 165.01 185.125 ;
      VIA 164.22 184.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 184.775 164.99 185.145 ;
      VIA 164.22 184.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 184.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 179.355 165.01 179.685 ;
      VIA 164.22 179.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 179.335 164.99 179.705 ;
      VIA 164.22 179.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 179.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 173.915 165.01 174.245 ;
      VIA 164.22 174.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 173.895 164.99 174.265 ;
      VIA 164.22 174.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 174.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 168.475 165.01 168.805 ;
      VIA 164.22 168.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 168.455 164.99 168.825 ;
      VIA 164.22 168.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 168.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 163.035 165.01 163.365 ;
      VIA 164.22 163.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 163.015 164.99 163.385 ;
      VIA 164.22 163.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 163.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 157.595 165.01 157.925 ;
      VIA 164.22 157.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 157.575 164.99 157.945 ;
      VIA 164.22 157.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 157.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 152.155 165.01 152.485 ;
      VIA 164.22 152.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 152.135 164.99 152.505 ;
      VIA 164.22 152.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 152.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 146.715 165.01 147.045 ;
      VIA 164.22 146.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 146.695 164.99 147.065 ;
      VIA 164.22 146.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 146.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 141.275 165.01 141.605 ;
      VIA 164.22 141.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 141.255 164.99 141.625 ;
      VIA 164.22 141.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 141.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 135.835 165.01 136.165 ;
      VIA 164.22 136 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 135.815 164.99 136.185 ;
      VIA 164.22 136 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 136 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 130.395 165.01 130.725 ;
      VIA 164.22 130.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 130.375 164.99 130.745 ;
      VIA 164.22 130.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 130.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 124.955 165.01 125.285 ;
      VIA 164.22 125.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 124.935 164.99 125.305 ;
      VIA 164.22 125.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 125.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 119.515 165.01 119.845 ;
      VIA 164.22 119.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 119.495 164.99 119.865 ;
      VIA 164.22 119.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 119.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 114.075 165.01 114.405 ;
      VIA 164.22 114.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 114.055 164.99 114.425 ;
      VIA 164.22 114.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 114.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 108.635 165.01 108.965 ;
      VIA 164.22 108.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 108.615 164.99 108.985 ;
      VIA 164.22 108.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 108.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 103.195 165.01 103.525 ;
      VIA 164.22 103.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 103.175 164.99 103.545 ;
      VIA 164.22 103.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 103.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 97.755 165.01 98.085 ;
      VIA 164.22 97.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 97.735 164.99 98.105 ;
      VIA 164.22 97.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 97.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 92.315 165.01 92.645 ;
      VIA 164.22 92.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 92.295 164.99 92.665 ;
      VIA 164.22 92.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 92.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 86.875 165.01 87.205 ;
      VIA 164.22 87.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 86.855 164.99 87.225 ;
      VIA 164.22 87.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 87.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 81.435 165.01 81.765 ;
      VIA 164.22 81.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 81.415 164.99 81.785 ;
      VIA 164.22 81.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 81.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 75.995 165.01 76.325 ;
      VIA 164.22 76.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 75.975 164.99 76.345 ;
      VIA 164.22 76.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 76.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 70.555 165.01 70.885 ;
      VIA 164.22 70.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 70.535 164.99 70.905 ;
      VIA 164.22 70.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 70.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 65.115 165.01 65.445 ;
      VIA 164.22 65.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 65.095 164.99 65.465 ;
      VIA 164.22 65.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 65.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 59.675 165.01 60.005 ;
      VIA 164.22 59.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 59.655 164.99 60.025 ;
      VIA 164.22 59.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 59.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 54.235 165.01 54.565 ;
      VIA 164.22 54.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 54.215 164.99 54.585 ;
      VIA 164.22 54.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 54.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 48.795 165.01 49.125 ;
      VIA 164.22 48.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 48.775 164.99 49.145 ;
      VIA 164.22 48.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 48.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 43.355 165.01 43.685 ;
      VIA 164.22 43.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 43.335 164.99 43.705 ;
      VIA 164.22 43.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 43.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 37.915 165.01 38.245 ;
      VIA 164.22 38.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 37.895 164.99 38.265 ;
      VIA 164.22 38.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 38.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 32.475 165.01 32.805 ;
      VIA 164.22 32.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 32.455 164.99 32.825 ;
      VIA 164.22 32.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 32.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 27.035 165.01 27.365 ;
      VIA 164.22 27.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 27.015 164.99 27.385 ;
      VIA 164.22 27.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 27.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 21.595 165.01 21.925 ;
      VIA 164.22 21.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 21.575 164.99 21.945 ;
      VIA 164.22 21.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 21.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 16.155 165.01 16.485 ;
      VIA 164.22 16.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 16.135 164.99 16.505 ;
      VIA 164.22 16.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 16.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 10.715 165.01 11.045 ;
      VIA 164.22 10.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 10.695 164.99 11.065 ;
      VIA 164.22 10.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 10.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  163.43 5.275 165.01 5.605 ;
      VIA 164.22 5.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  163.45 5.255 164.99 5.625 ;
      VIA 164.22 5.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 164.22 5.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 701.595 137.87 701.925 ;
      VIA 137.08 701.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 701.575 137.85 701.945 ;
      VIA 137.08 701.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 701.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 696.155 137.87 696.485 ;
      VIA 137.08 696.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 696.135 137.85 696.505 ;
      VIA 137.08 696.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 696.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 690.715 137.87 691.045 ;
      VIA 137.08 690.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 690.695 137.85 691.065 ;
      VIA 137.08 690.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 690.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 685.275 137.87 685.605 ;
      VIA 137.08 685.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 685.255 137.85 685.625 ;
      VIA 137.08 685.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 685.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 679.835 137.87 680.165 ;
      VIA 137.08 680 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 679.815 137.85 680.185 ;
      VIA 137.08 680 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 680 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 674.395 137.87 674.725 ;
      VIA 137.08 674.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 674.375 137.85 674.745 ;
      VIA 137.08 674.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 674.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 668.955 137.87 669.285 ;
      VIA 137.08 669.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 668.935 137.85 669.305 ;
      VIA 137.08 669.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 669.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 663.515 137.87 663.845 ;
      VIA 137.08 663.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 663.495 137.85 663.865 ;
      VIA 137.08 663.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 663.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 658.075 137.87 658.405 ;
      VIA 137.08 658.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 658.055 137.85 658.425 ;
      VIA 137.08 658.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 658.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 652.635 137.87 652.965 ;
      VIA 137.08 652.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 652.615 137.85 652.985 ;
      VIA 137.08 652.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 652.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 647.195 137.87 647.525 ;
      VIA 137.08 647.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 647.175 137.85 647.545 ;
      VIA 137.08 647.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 647.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 641.755 137.87 642.085 ;
      VIA 137.08 641.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 641.735 137.85 642.105 ;
      VIA 137.08 641.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 641.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 636.315 137.87 636.645 ;
      VIA 137.08 636.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 636.295 137.85 636.665 ;
      VIA 137.08 636.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 636.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 630.875 137.87 631.205 ;
      VIA 137.08 631.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 630.855 137.85 631.225 ;
      VIA 137.08 631.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 631.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 625.435 137.87 625.765 ;
      VIA 137.08 625.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 625.415 137.85 625.785 ;
      VIA 137.08 625.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 625.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 619.995 137.87 620.325 ;
      VIA 137.08 620.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 619.975 137.85 620.345 ;
      VIA 137.08 620.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 620.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 614.555 137.87 614.885 ;
      VIA 137.08 614.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 614.535 137.85 614.905 ;
      VIA 137.08 614.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 614.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 609.115 137.87 609.445 ;
      VIA 137.08 609.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 609.095 137.85 609.465 ;
      VIA 137.08 609.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 609.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 603.675 137.87 604.005 ;
      VIA 137.08 603.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 603.655 137.85 604.025 ;
      VIA 137.08 603.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 603.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 598.235 137.87 598.565 ;
      VIA 137.08 598.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 598.215 137.85 598.585 ;
      VIA 137.08 598.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 598.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 592.795 137.87 593.125 ;
      VIA 137.08 592.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 592.775 137.85 593.145 ;
      VIA 137.08 592.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 592.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 587.355 137.87 587.685 ;
      VIA 137.08 587.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 587.335 137.85 587.705 ;
      VIA 137.08 587.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 587.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 581.915 137.87 582.245 ;
      VIA 137.08 582.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 581.895 137.85 582.265 ;
      VIA 137.08 582.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 582.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 576.475 137.87 576.805 ;
      VIA 137.08 576.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 576.455 137.85 576.825 ;
      VIA 137.08 576.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 576.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 571.035 137.87 571.365 ;
      VIA 137.08 571.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 571.015 137.85 571.385 ;
      VIA 137.08 571.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 571.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 565.595 137.87 565.925 ;
      VIA 137.08 565.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 565.575 137.85 565.945 ;
      VIA 137.08 565.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 565.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 560.155 137.87 560.485 ;
      VIA 137.08 560.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 560.135 137.85 560.505 ;
      VIA 137.08 560.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 560.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 554.715 137.87 555.045 ;
      VIA 137.08 554.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 554.695 137.85 555.065 ;
      VIA 137.08 554.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 554.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 549.275 137.87 549.605 ;
      VIA 137.08 549.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 549.255 137.85 549.625 ;
      VIA 137.08 549.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 549.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 543.835 137.87 544.165 ;
      VIA 137.08 544 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 543.815 137.85 544.185 ;
      VIA 137.08 544 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 544 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 538.395 137.87 538.725 ;
      VIA 137.08 538.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 538.375 137.85 538.745 ;
      VIA 137.08 538.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 538.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 532.955 137.87 533.285 ;
      VIA 137.08 533.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 532.935 137.85 533.305 ;
      VIA 137.08 533.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 533.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 527.515 137.87 527.845 ;
      VIA 137.08 527.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 527.495 137.85 527.865 ;
      VIA 137.08 527.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 527.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 522.075 137.87 522.405 ;
      VIA 137.08 522.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 522.055 137.85 522.425 ;
      VIA 137.08 522.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 522.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 516.635 137.87 516.965 ;
      VIA 137.08 516.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 516.615 137.85 516.985 ;
      VIA 137.08 516.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 516.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 511.195 137.87 511.525 ;
      VIA 137.08 511.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 511.175 137.85 511.545 ;
      VIA 137.08 511.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 511.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 505.755 137.87 506.085 ;
      VIA 137.08 505.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 505.735 137.85 506.105 ;
      VIA 137.08 505.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 505.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 500.315 137.87 500.645 ;
      VIA 137.08 500.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 500.295 137.85 500.665 ;
      VIA 137.08 500.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 500.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 494.875 137.87 495.205 ;
      VIA 137.08 495.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 494.855 137.85 495.225 ;
      VIA 137.08 495.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 495.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 489.435 137.87 489.765 ;
      VIA 137.08 489.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 489.415 137.85 489.785 ;
      VIA 137.08 489.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 489.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 483.995 137.87 484.325 ;
      VIA 137.08 484.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 483.975 137.85 484.345 ;
      VIA 137.08 484.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 484.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 478.555 137.87 478.885 ;
      VIA 137.08 478.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 478.535 137.85 478.905 ;
      VIA 137.08 478.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 478.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 473.115 137.87 473.445 ;
      VIA 137.08 473.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 473.095 137.85 473.465 ;
      VIA 137.08 473.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 473.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 467.675 137.87 468.005 ;
      VIA 137.08 467.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 467.655 137.85 468.025 ;
      VIA 137.08 467.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 467.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 462.235 137.87 462.565 ;
      VIA 137.08 462.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 462.215 137.85 462.585 ;
      VIA 137.08 462.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 462.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 456.795 137.87 457.125 ;
      VIA 137.08 456.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 456.775 137.85 457.145 ;
      VIA 137.08 456.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 456.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 451.355 137.87 451.685 ;
      VIA 137.08 451.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 451.335 137.85 451.705 ;
      VIA 137.08 451.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 451.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 445.915 137.87 446.245 ;
      VIA 137.08 446.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 445.895 137.85 446.265 ;
      VIA 137.08 446.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 446.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 440.475 137.87 440.805 ;
      VIA 137.08 440.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 440.455 137.85 440.825 ;
      VIA 137.08 440.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 440.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 435.035 137.87 435.365 ;
      VIA 137.08 435.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 435.015 137.85 435.385 ;
      VIA 137.08 435.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 435.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 429.595 137.87 429.925 ;
      VIA 137.08 429.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 429.575 137.85 429.945 ;
      VIA 137.08 429.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 429.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 424.155 137.87 424.485 ;
      VIA 137.08 424.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 424.135 137.85 424.505 ;
      VIA 137.08 424.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 424.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 418.715 137.87 419.045 ;
      VIA 137.08 418.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 418.695 137.85 419.065 ;
      VIA 137.08 418.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 418.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 413.275 137.87 413.605 ;
      VIA 137.08 413.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 413.255 137.85 413.625 ;
      VIA 137.08 413.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 413.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 407.835 137.87 408.165 ;
      VIA 137.08 408 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 407.815 137.85 408.185 ;
      VIA 137.08 408 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 408 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 402.395 137.87 402.725 ;
      VIA 137.08 402.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 402.375 137.85 402.745 ;
      VIA 137.08 402.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 402.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 396.955 137.87 397.285 ;
      VIA 137.08 397.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 396.935 137.85 397.305 ;
      VIA 137.08 397.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 397.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 391.515 137.87 391.845 ;
      VIA 137.08 391.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 391.495 137.85 391.865 ;
      VIA 137.08 391.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 391.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 386.075 137.87 386.405 ;
      VIA 137.08 386.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 386.055 137.85 386.425 ;
      VIA 137.08 386.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 386.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 380.635 137.87 380.965 ;
      VIA 137.08 380.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 380.615 137.85 380.985 ;
      VIA 137.08 380.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 380.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 375.195 137.87 375.525 ;
      VIA 137.08 375.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 375.175 137.85 375.545 ;
      VIA 137.08 375.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 375.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 369.755 137.87 370.085 ;
      VIA 137.08 369.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 369.735 137.85 370.105 ;
      VIA 137.08 369.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 369.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 364.315 137.87 364.645 ;
      VIA 137.08 364.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 364.295 137.85 364.665 ;
      VIA 137.08 364.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 364.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 358.875 137.87 359.205 ;
      VIA 137.08 359.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 358.855 137.85 359.225 ;
      VIA 137.08 359.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 359.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 353.435 137.87 353.765 ;
      VIA 137.08 353.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 353.415 137.85 353.785 ;
      VIA 137.08 353.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 353.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 347.995 137.87 348.325 ;
      VIA 137.08 348.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 347.975 137.85 348.345 ;
      VIA 137.08 348.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 348.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 342.555 137.87 342.885 ;
      VIA 137.08 342.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 342.535 137.85 342.905 ;
      VIA 137.08 342.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 342.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 337.115 137.87 337.445 ;
      VIA 137.08 337.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 337.095 137.85 337.465 ;
      VIA 137.08 337.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 337.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 331.675 137.87 332.005 ;
      VIA 137.08 331.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 331.655 137.85 332.025 ;
      VIA 137.08 331.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 331.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 326.235 137.87 326.565 ;
      VIA 137.08 326.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 326.215 137.85 326.585 ;
      VIA 137.08 326.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 326.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 320.795 137.87 321.125 ;
      VIA 137.08 320.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 320.775 137.85 321.145 ;
      VIA 137.08 320.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 320.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 315.355 137.87 315.685 ;
      VIA 137.08 315.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 315.335 137.85 315.705 ;
      VIA 137.08 315.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 315.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 309.915 137.87 310.245 ;
      VIA 137.08 310.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 309.895 137.85 310.265 ;
      VIA 137.08 310.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 310.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 304.475 137.87 304.805 ;
      VIA 137.08 304.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 304.455 137.85 304.825 ;
      VIA 137.08 304.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 304.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 299.035 137.87 299.365 ;
      VIA 137.08 299.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 299.015 137.85 299.385 ;
      VIA 137.08 299.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 299.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 293.595 137.87 293.925 ;
      VIA 137.08 293.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 293.575 137.85 293.945 ;
      VIA 137.08 293.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 293.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 288.155 137.87 288.485 ;
      VIA 137.08 288.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 288.135 137.85 288.505 ;
      VIA 137.08 288.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 288.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 282.715 137.87 283.045 ;
      VIA 137.08 282.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 282.695 137.85 283.065 ;
      VIA 137.08 282.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 282.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 277.275 137.87 277.605 ;
      VIA 137.08 277.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 277.255 137.85 277.625 ;
      VIA 137.08 277.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 277.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 271.835 137.87 272.165 ;
      VIA 137.08 272 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 271.815 137.85 272.185 ;
      VIA 137.08 272 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 272 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 266.395 137.87 266.725 ;
      VIA 137.08 266.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 266.375 137.85 266.745 ;
      VIA 137.08 266.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 266.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 260.955 137.87 261.285 ;
      VIA 137.08 261.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 260.935 137.85 261.305 ;
      VIA 137.08 261.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 261.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 255.515 137.87 255.845 ;
      VIA 137.08 255.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 255.495 137.85 255.865 ;
      VIA 137.08 255.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 255.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 250.075 137.87 250.405 ;
      VIA 137.08 250.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 250.055 137.85 250.425 ;
      VIA 137.08 250.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 250.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 244.635 137.87 244.965 ;
      VIA 137.08 244.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 244.615 137.85 244.985 ;
      VIA 137.08 244.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 244.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 239.195 137.87 239.525 ;
      VIA 137.08 239.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 239.175 137.85 239.545 ;
      VIA 137.08 239.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 239.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 233.755 137.87 234.085 ;
      VIA 137.08 233.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 233.735 137.85 234.105 ;
      VIA 137.08 233.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 233.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 228.315 137.87 228.645 ;
      VIA 137.08 228.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 228.295 137.85 228.665 ;
      VIA 137.08 228.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 228.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 222.875 137.87 223.205 ;
      VIA 137.08 223.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 222.855 137.85 223.225 ;
      VIA 137.08 223.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 223.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 217.435 137.87 217.765 ;
      VIA 137.08 217.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 217.415 137.85 217.785 ;
      VIA 137.08 217.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 217.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 211.995 137.87 212.325 ;
      VIA 137.08 212.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 211.975 137.85 212.345 ;
      VIA 137.08 212.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 212.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 206.555 137.87 206.885 ;
      VIA 137.08 206.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 206.535 137.85 206.905 ;
      VIA 137.08 206.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 206.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 201.115 137.87 201.445 ;
      VIA 137.08 201.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 201.095 137.85 201.465 ;
      VIA 137.08 201.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 201.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 195.675 137.87 196.005 ;
      VIA 137.08 195.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 195.655 137.85 196.025 ;
      VIA 137.08 195.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 195.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 190.235 137.87 190.565 ;
      VIA 137.08 190.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 190.215 137.85 190.585 ;
      VIA 137.08 190.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 190.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 184.795 137.87 185.125 ;
      VIA 137.08 184.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 184.775 137.85 185.145 ;
      VIA 137.08 184.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 184.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 179.355 137.87 179.685 ;
      VIA 137.08 179.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 179.335 137.85 179.705 ;
      VIA 137.08 179.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 179.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 173.915 137.87 174.245 ;
      VIA 137.08 174.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 173.895 137.85 174.265 ;
      VIA 137.08 174.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 174.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 168.475 137.87 168.805 ;
      VIA 137.08 168.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 168.455 137.85 168.825 ;
      VIA 137.08 168.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 168.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 163.035 137.87 163.365 ;
      VIA 137.08 163.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 163.015 137.85 163.385 ;
      VIA 137.08 163.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 163.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 157.595 137.87 157.925 ;
      VIA 137.08 157.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 157.575 137.85 157.945 ;
      VIA 137.08 157.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 157.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 152.155 137.87 152.485 ;
      VIA 137.08 152.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 152.135 137.85 152.505 ;
      VIA 137.08 152.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 152.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 146.715 137.87 147.045 ;
      VIA 137.08 146.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 146.695 137.85 147.065 ;
      VIA 137.08 146.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 146.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 141.275 137.87 141.605 ;
      VIA 137.08 141.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 141.255 137.85 141.625 ;
      VIA 137.08 141.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 141.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 135.835 137.87 136.165 ;
      VIA 137.08 136 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 135.815 137.85 136.185 ;
      VIA 137.08 136 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 136 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 130.395 137.87 130.725 ;
      VIA 137.08 130.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 130.375 137.85 130.745 ;
      VIA 137.08 130.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 130.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 124.955 137.87 125.285 ;
      VIA 137.08 125.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 124.935 137.85 125.305 ;
      VIA 137.08 125.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 125.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 119.515 137.87 119.845 ;
      VIA 137.08 119.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 119.495 137.85 119.865 ;
      VIA 137.08 119.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 119.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 114.075 137.87 114.405 ;
      VIA 137.08 114.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 114.055 137.85 114.425 ;
      VIA 137.08 114.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 114.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 108.635 137.87 108.965 ;
      VIA 137.08 108.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 108.615 137.85 108.985 ;
      VIA 137.08 108.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 108.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 103.195 137.87 103.525 ;
      VIA 137.08 103.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 103.175 137.85 103.545 ;
      VIA 137.08 103.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 103.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 97.755 137.87 98.085 ;
      VIA 137.08 97.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 97.735 137.85 98.105 ;
      VIA 137.08 97.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 97.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 92.315 137.87 92.645 ;
      VIA 137.08 92.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 92.295 137.85 92.665 ;
      VIA 137.08 92.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 92.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 86.875 137.87 87.205 ;
      VIA 137.08 87.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 86.855 137.85 87.225 ;
      VIA 137.08 87.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 87.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 81.435 137.87 81.765 ;
      VIA 137.08 81.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 81.415 137.85 81.785 ;
      VIA 137.08 81.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 81.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 75.995 137.87 76.325 ;
      VIA 137.08 76.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 75.975 137.85 76.345 ;
      VIA 137.08 76.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 76.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 70.555 137.87 70.885 ;
      VIA 137.08 70.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 70.535 137.85 70.905 ;
      VIA 137.08 70.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 70.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 65.115 137.87 65.445 ;
      VIA 137.08 65.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 65.095 137.85 65.465 ;
      VIA 137.08 65.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 65.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 59.675 137.87 60.005 ;
      VIA 137.08 59.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 59.655 137.85 60.025 ;
      VIA 137.08 59.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 59.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 54.235 137.87 54.565 ;
      VIA 137.08 54.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 54.215 137.85 54.585 ;
      VIA 137.08 54.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 54.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 48.795 137.87 49.125 ;
      VIA 137.08 48.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 48.775 137.85 49.145 ;
      VIA 137.08 48.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 48.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 43.355 137.87 43.685 ;
      VIA 137.08 43.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 43.335 137.85 43.705 ;
      VIA 137.08 43.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 43.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 37.915 137.87 38.245 ;
      VIA 137.08 38.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 37.895 137.85 38.265 ;
      VIA 137.08 38.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 38.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 32.475 137.87 32.805 ;
      VIA 137.08 32.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 32.455 137.85 32.825 ;
      VIA 137.08 32.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 32.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 27.035 137.87 27.365 ;
      VIA 137.08 27.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 27.015 137.85 27.385 ;
      VIA 137.08 27.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 27.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 21.595 137.87 21.925 ;
      VIA 137.08 21.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 21.575 137.85 21.945 ;
      VIA 137.08 21.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 21.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 16.155 137.87 16.485 ;
      VIA 137.08 16.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 16.135 137.85 16.505 ;
      VIA 137.08 16.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 16.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 10.715 137.87 11.045 ;
      VIA 137.08 10.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 10.695 137.85 11.065 ;
      VIA 137.08 10.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 10.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  136.29 5.275 137.87 5.605 ;
      VIA 137.08 5.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  136.31 5.255 137.85 5.625 ;
      VIA 137.08 5.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 137.08 5.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 701.595 110.73 701.925 ;
      VIA 109.94 701.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 701.575 110.71 701.945 ;
      VIA 109.94 701.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 701.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 696.155 110.73 696.485 ;
      VIA 109.94 696.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 696.135 110.71 696.505 ;
      VIA 109.94 696.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 696.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 690.715 110.73 691.045 ;
      VIA 109.94 690.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 690.695 110.71 691.065 ;
      VIA 109.94 690.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 690.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 685.275 110.73 685.605 ;
      VIA 109.94 685.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 685.255 110.71 685.625 ;
      VIA 109.94 685.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 685.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 679.835 110.73 680.165 ;
      VIA 109.94 680 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 679.815 110.71 680.185 ;
      VIA 109.94 680 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 680 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 674.395 110.73 674.725 ;
      VIA 109.94 674.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 674.375 110.71 674.745 ;
      VIA 109.94 674.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 674.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 668.955 110.73 669.285 ;
      VIA 109.94 669.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 668.935 110.71 669.305 ;
      VIA 109.94 669.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 669.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 663.515 110.73 663.845 ;
      VIA 109.94 663.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 663.495 110.71 663.865 ;
      VIA 109.94 663.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 663.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 658.075 110.73 658.405 ;
      VIA 109.94 658.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 658.055 110.71 658.425 ;
      VIA 109.94 658.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 658.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 652.635 110.73 652.965 ;
      VIA 109.94 652.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 652.615 110.71 652.985 ;
      VIA 109.94 652.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 652.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 647.195 110.73 647.525 ;
      VIA 109.94 647.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 647.175 110.71 647.545 ;
      VIA 109.94 647.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 647.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 641.755 110.73 642.085 ;
      VIA 109.94 641.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 641.735 110.71 642.105 ;
      VIA 109.94 641.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 641.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 636.315 110.73 636.645 ;
      VIA 109.94 636.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 636.295 110.71 636.665 ;
      VIA 109.94 636.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 636.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 630.875 110.73 631.205 ;
      VIA 109.94 631.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 630.855 110.71 631.225 ;
      VIA 109.94 631.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 631.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 625.435 110.73 625.765 ;
      VIA 109.94 625.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 625.415 110.71 625.785 ;
      VIA 109.94 625.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 625.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 619.995 110.73 620.325 ;
      VIA 109.94 620.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 619.975 110.71 620.345 ;
      VIA 109.94 620.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 620.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 614.555 110.73 614.885 ;
      VIA 109.94 614.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 614.535 110.71 614.905 ;
      VIA 109.94 614.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 614.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 609.115 110.73 609.445 ;
      VIA 109.94 609.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 609.095 110.71 609.465 ;
      VIA 109.94 609.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 609.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 603.675 110.73 604.005 ;
      VIA 109.94 603.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 603.655 110.71 604.025 ;
      VIA 109.94 603.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 603.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 598.235 110.73 598.565 ;
      VIA 109.94 598.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 598.215 110.71 598.585 ;
      VIA 109.94 598.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 598.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 592.795 110.73 593.125 ;
      VIA 109.94 592.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 592.775 110.71 593.145 ;
      VIA 109.94 592.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 592.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 587.355 110.73 587.685 ;
      VIA 109.94 587.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 587.335 110.71 587.705 ;
      VIA 109.94 587.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 587.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 581.915 110.73 582.245 ;
      VIA 109.94 582.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 581.895 110.71 582.265 ;
      VIA 109.94 582.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 582.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 576.475 110.73 576.805 ;
      VIA 109.94 576.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 576.455 110.71 576.825 ;
      VIA 109.94 576.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 576.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 571.035 110.73 571.365 ;
      VIA 109.94 571.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 571.015 110.71 571.385 ;
      VIA 109.94 571.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 571.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 565.595 110.73 565.925 ;
      VIA 109.94 565.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 565.575 110.71 565.945 ;
      VIA 109.94 565.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 565.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 560.155 110.73 560.485 ;
      VIA 109.94 560.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 560.135 110.71 560.505 ;
      VIA 109.94 560.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 560.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 554.715 110.73 555.045 ;
      VIA 109.94 554.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 554.695 110.71 555.065 ;
      VIA 109.94 554.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 554.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 549.275 110.73 549.605 ;
      VIA 109.94 549.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 549.255 110.71 549.625 ;
      VIA 109.94 549.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 549.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 543.835 110.73 544.165 ;
      VIA 109.94 544 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 543.815 110.71 544.185 ;
      VIA 109.94 544 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 544 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 538.395 110.73 538.725 ;
      VIA 109.94 538.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 538.375 110.71 538.745 ;
      VIA 109.94 538.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 538.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 532.955 110.73 533.285 ;
      VIA 109.94 533.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 532.935 110.71 533.305 ;
      VIA 109.94 533.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 533.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 527.515 110.73 527.845 ;
      VIA 109.94 527.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 527.495 110.71 527.865 ;
      VIA 109.94 527.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 527.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 522.075 110.73 522.405 ;
      VIA 109.94 522.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 522.055 110.71 522.425 ;
      VIA 109.94 522.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 522.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 516.635 110.73 516.965 ;
      VIA 109.94 516.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 516.615 110.71 516.985 ;
      VIA 109.94 516.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 516.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 511.195 110.73 511.525 ;
      VIA 109.94 511.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 511.175 110.71 511.545 ;
      VIA 109.94 511.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 511.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 505.755 110.73 506.085 ;
      VIA 109.94 505.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 505.735 110.71 506.105 ;
      VIA 109.94 505.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 505.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 500.315 110.73 500.645 ;
      VIA 109.94 500.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 500.295 110.71 500.665 ;
      VIA 109.94 500.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 500.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 494.875 110.73 495.205 ;
      VIA 109.94 495.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 494.855 110.71 495.225 ;
      VIA 109.94 495.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 495.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 489.435 110.73 489.765 ;
      VIA 109.94 489.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 489.415 110.71 489.785 ;
      VIA 109.94 489.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 489.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 483.995 110.73 484.325 ;
      VIA 109.94 484.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 483.975 110.71 484.345 ;
      VIA 109.94 484.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 484.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 478.555 110.73 478.885 ;
      VIA 109.94 478.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 478.535 110.71 478.905 ;
      VIA 109.94 478.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 478.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 473.115 110.73 473.445 ;
      VIA 109.94 473.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 473.095 110.71 473.465 ;
      VIA 109.94 473.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 473.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 467.675 110.73 468.005 ;
      VIA 109.94 467.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 467.655 110.71 468.025 ;
      VIA 109.94 467.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 467.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 462.235 110.73 462.565 ;
      VIA 109.94 462.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 462.215 110.71 462.585 ;
      VIA 109.94 462.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 462.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 456.795 110.73 457.125 ;
      VIA 109.94 456.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 456.775 110.71 457.145 ;
      VIA 109.94 456.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 456.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 451.355 110.73 451.685 ;
      VIA 109.94 451.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 451.335 110.71 451.705 ;
      VIA 109.94 451.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 451.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 445.915 110.73 446.245 ;
      VIA 109.94 446.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 445.895 110.71 446.265 ;
      VIA 109.94 446.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 446.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 440.475 110.73 440.805 ;
      VIA 109.94 440.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 440.455 110.71 440.825 ;
      VIA 109.94 440.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 440.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 435.035 110.73 435.365 ;
      VIA 109.94 435.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 435.015 110.71 435.385 ;
      VIA 109.94 435.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 435.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 429.595 110.73 429.925 ;
      VIA 109.94 429.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 429.575 110.71 429.945 ;
      VIA 109.94 429.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 429.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 424.155 110.73 424.485 ;
      VIA 109.94 424.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 424.135 110.71 424.505 ;
      VIA 109.94 424.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 424.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 418.715 110.73 419.045 ;
      VIA 109.94 418.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 418.695 110.71 419.065 ;
      VIA 109.94 418.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 418.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 413.275 110.73 413.605 ;
      VIA 109.94 413.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 413.255 110.71 413.625 ;
      VIA 109.94 413.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 413.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 407.835 110.73 408.165 ;
      VIA 109.94 408 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 407.815 110.71 408.185 ;
      VIA 109.94 408 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 408 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 402.395 110.73 402.725 ;
      VIA 109.94 402.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 402.375 110.71 402.745 ;
      VIA 109.94 402.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 402.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 396.955 110.73 397.285 ;
      VIA 109.94 397.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 396.935 110.71 397.305 ;
      VIA 109.94 397.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 397.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 391.515 110.73 391.845 ;
      VIA 109.94 391.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 391.495 110.71 391.865 ;
      VIA 109.94 391.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 391.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 386.075 110.73 386.405 ;
      VIA 109.94 386.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 386.055 110.71 386.425 ;
      VIA 109.94 386.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 386.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 380.635 110.73 380.965 ;
      VIA 109.94 380.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 380.615 110.71 380.985 ;
      VIA 109.94 380.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 380.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 375.195 110.73 375.525 ;
      VIA 109.94 375.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 375.175 110.71 375.545 ;
      VIA 109.94 375.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 375.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 369.755 110.73 370.085 ;
      VIA 109.94 369.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 369.735 110.71 370.105 ;
      VIA 109.94 369.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 369.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 364.315 110.73 364.645 ;
      VIA 109.94 364.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 364.295 110.71 364.665 ;
      VIA 109.94 364.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 364.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 358.875 110.73 359.205 ;
      VIA 109.94 359.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 358.855 110.71 359.225 ;
      VIA 109.94 359.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 359.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 353.435 110.73 353.765 ;
      VIA 109.94 353.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 353.415 110.71 353.785 ;
      VIA 109.94 353.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 353.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 347.995 110.73 348.325 ;
      VIA 109.94 348.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 347.975 110.71 348.345 ;
      VIA 109.94 348.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 348.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 342.555 110.73 342.885 ;
      VIA 109.94 342.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 342.535 110.71 342.905 ;
      VIA 109.94 342.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 342.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 337.115 110.73 337.445 ;
      VIA 109.94 337.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 337.095 110.71 337.465 ;
      VIA 109.94 337.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 337.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 331.675 110.73 332.005 ;
      VIA 109.94 331.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 331.655 110.71 332.025 ;
      VIA 109.94 331.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 331.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 326.235 110.73 326.565 ;
      VIA 109.94 326.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 326.215 110.71 326.585 ;
      VIA 109.94 326.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 326.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 320.795 110.73 321.125 ;
      VIA 109.94 320.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 320.775 110.71 321.145 ;
      VIA 109.94 320.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 320.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 315.355 110.73 315.685 ;
      VIA 109.94 315.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 315.335 110.71 315.705 ;
      VIA 109.94 315.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 315.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 309.915 110.73 310.245 ;
      VIA 109.94 310.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 309.895 110.71 310.265 ;
      VIA 109.94 310.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 310.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 304.475 110.73 304.805 ;
      VIA 109.94 304.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 304.455 110.71 304.825 ;
      VIA 109.94 304.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 304.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 299.035 110.73 299.365 ;
      VIA 109.94 299.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 299.015 110.71 299.385 ;
      VIA 109.94 299.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 299.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 293.595 110.73 293.925 ;
      VIA 109.94 293.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 293.575 110.71 293.945 ;
      VIA 109.94 293.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 293.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 288.155 110.73 288.485 ;
      VIA 109.94 288.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 288.135 110.71 288.505 ;
      VIA 109.94 288.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 288.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 282.715 110.73 283.045 ;
      VIA 109.94 282.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 282.695 110.71 283.065 ;
      VIA 109.94 282.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 282.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 277.275 110.73 277.605 ;
      VIA 109.94 277.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 277.255 110.71 277.625 ;
      VIA 109.94 277.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 277.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 271.835 110.73 272.165 ;
      VIA 109.94 272 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 271.815 110.71 272.185 ;
      VIA 109.94 272 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 272 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 266.395 110.73 266.725 ;
      VIA 109.94 266.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 266.375 110.71 266.745 ;
      VIA 109.94 266.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 266.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 260.955 110.73 261.285 ;
      VIA 109.94 261.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 260.935 110.71 261.305 ;
      VIA 109.94 261.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 261.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 255.515 110.73 255.845 ;
      VIA 109.94 255.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 255.495 110.71 255.865 ;
      VIA 109.94 255.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 255.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 250.075 110.73 250.405 ;
      VIA 109.94 250.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 250.055 110.71 250.425 ;
      VIA 109.94 250.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 250.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 244.635 110.73 244.965 ;
      VIA 109.94 244.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 244.615 110.71 244.985 ;
      VIA 109.94 244.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 244.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 239.195 110.73 239.525 ;
      VIA 109.94 239.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 239.175 110.71 239.545 ;
      VIA 109.94 239.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 239.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 233.755 110.73 234.085 ;
      VIA 109.94 233.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 233.735 110.71 234.105 ;
      VIA 109.94 233.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 233.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 228.315 110.73 228.645 ;
      VIA 109.94 228.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 228.295 110.71 228.665 ;
      VIA 109.94 228.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 228.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 222.875 110.73 223.205 ;
      VIA 109.94 223.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 222.855 110.71 223.225 ;
      VIA 109.94 223.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 223.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 217.435 110.73 217.765 ;
      VIA 109.94 217.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 217.415 110.71 217.785 ;
      VIA 109.94 217.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 217.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 211.995 110.73 212.325 ;
      VIA 109.94 212.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 211.975 110.71 212.345 ;
      VIA 109.94 212.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 212.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 206.555 110.73 206.885 ;
      VIA 109.94 206.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 206.535 110.71 206.905 ;
      VIA 109.94 206.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 206.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 201.115 110.73 201.445 ;
      VIA 109.94 201.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 201.095 110.71 201.465 ;
      VIA 109.94 201.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 201.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 195.675 110.73 196.005 ;
      VIA 109.94 195.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 195.655 110.71 196.025 ;
      VIA 109.94 195.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 195.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 190.235 110.73 190.565 ;
      VIA 109.94 190.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 190.215 110.71 190.585 ;
      VIA 109.94 190.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 190.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 184.795 110.73 185.125 ;
      VIA 109.94 184.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 184.775 110.71 185.145 ;
      VIA 109.94 184.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 184.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 179.355 110.73 179.685 ;
      VIA 109.94 179.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 179.335 110.71 179.705 ;
      VIA 109.94 179.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 179.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 173.915 110.73 174.245 ;
      VIA 109.94 174.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 173.895 110.71 174.265 ;
      VIA 109.94 174.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 174.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 168.475 110.73 168.805 ;
      VIA 109.94 168.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 168.455 110.71 168.825 ;
      VIA 109.94 168.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 168.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 163.035 110.73 163.365 ;
      VIA 109.94 163.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 163.015 110.71 163.385 ;
      VIA 109.94 163.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 163.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 157.595 110.73 157.925 ;
      VIA 109.94 157.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 157.575 110.71 157.945 ;
      VIA 109.94 157.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 157.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 152.155 110.73 152.485 ;
      VIA 109.94 152.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 152.135 110.71 152.505 ;
      VIA 109.94 152.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 152.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 146.715 110.73 147.045 ;
      VIA 109.94 146.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 146.695 110.71 147.065 ;
      VIA 109.94 146.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 146.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 141.275 110.73 141.605 ;
      VIA 109.94 141.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 141.255 110.71 141.625 ;
      VIA 109.94 141.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 141.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 135.835 110.73 136.165 ;
      VIA 109.94 136 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 135.815 110.71 136.185 ;
      VIA 109.94 136 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 136 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 130.395 110.73 130.725 ;
      VIA 109.94 130.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 130.375 110.71 130.745 ;
      VIA 109.94 130.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 130.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 124.955 110.73 125.285 ;
      VIA 109.94 125.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 124.935 110.71 125.305 ;
      VIA 109.94 125.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 125.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 119.515 110.73 119.845 ;
      VIA 109.94 119.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 119.495 110.71 119.865 ;
      VIA 109.94 119.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 119.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 114.075 110.73 114.405 ;
      VIA 109.94 114.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 114.055 110.71 114.425 ;
      VIA 109.94 114.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 114.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 108.635 110.73 108.965 ;
      VIA 109.94 108.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 108.615 110.71 108.985 ;
      VIA 109.94 108.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 108.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 103.195 110.73 103.525 ;
      VIA 109.94 103.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 103.175 110.71 103.545 ;
      VIA 109.94 103.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 103.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 97.755 110.73 98.085 ;
      VIA 109.94 97.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 97.735 110.71 98.105 ;
      VIA 109.94 97.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 97.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 92.315 110.73 92.645 ;
      VIA 109.94 92.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 92.295 110.71 92.665 ;
      VIA 109.94 92.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 92.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 86.875 110.73 87.205 ;
      VIA 109.94 87.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 86.855 110.71 87.225 ;
      VIA 109.94 87.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 87.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 81.435 110.73 81.765 ;
      VIA 109.94 81.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 81.415 110.71 81.785 ;
      VIA 109.94 81.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 81.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 75.995 110.73 76.325 ;
      VIA 109.94 76.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 75.975 110.71 76.345 ;
      VIA 109.94 76.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 76.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 70.555 110.73 70.885 ;
      VIA 109.94 70.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 70.535 110.71 70.905 ;
      VIA 109.94 70.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 70.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 65.115 110.73 65.445 ;
      VIA 109.94 65.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 65.095 110.71 65.465 ;
      VIA 109.94 65.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 65.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 59.675 110.73 60.005 ;
      VIA 109.94 59.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 59.655 110.71 60.025 ;
      VIA 109.94 59.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 59.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 54.235 110.73 54.565 ;
      VIA 109.94 54.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 54.215 110.71 54.585 ;
      VIA 109.94 54.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 54.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 48.795 110.73 49.125 ;
      VIA 109.94 48.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 48.775 110.71 49.145 ;
      VIA 109.94 48.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 48.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 43.355 110.73 43.685 ;
      VIA 109.94 43.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 43.335 110.71 43.705 ;
      VIA 109.94 43.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 43.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 37.915 110.73 38.245 ;
      VIA 109.94 38.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 37.895 110.71 38.265 ;
      VIA 109.94 38.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 38.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 32.475 110.73 32.805 ;
      VIA 109.94 32.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 32.455 110.71 32.825 ;
      VIA 109.94 32.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 32.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 27.035 110.73 27.365 ;
      VIA 109.94 27.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 27.015 110.71 27.385 ;
      VIA 109.94 27.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 27.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 21.595 110.73 21.925 ;
      VIA 109.94 21.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 21.575 110.71 21.945 ;
      VIA 109.94 21.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 21.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 16.155 110.73 16.485 ;
      VIA 109.94 16.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 16.135 110.71 16.505 ;
      VIA 109.94 16.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 16.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 10.715 110.73 11.045 ;
      VIA 109.94 10.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 10.695 110.71 11.065 ;
      VIA 109.94 10.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 10.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  109.15 5.275 110.73 5.605 ;
      VIA 109.94 5.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  109.17 5.255 110.71 5.625 ;
      VIA 109.94 5.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 109.94 5.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 701.595 83.59 701.925 ;
      VIA 82.8 701.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 701.575 83.57 701.945 ;
      VIA 82.8 701.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 701.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 696.155 83.59 696.485 ;
      VIA 82.8 696.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 696.135 83.57 696.505 ;
      VIA 82.8 696.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 696.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 690.715 83.59 691.045 ;
      VIA 82.8 690.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 690.695 83.57 691.065 ;
      VIA 82.8 690.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 690.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 685.275 83.59 685.605 ;
      VIA 82.8 685.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 685.255 83.57 685.625 ;
      VIA 82.8 685.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 685.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 679.835 83.59 680.165 ;
      VIA 82.8 680 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 679.815 83.57 680.185 ;
      VIA 82.8 680 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 680 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 674.395 83.59 674.725 ;
      VIA 82.8 674.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 674.375 83.57 674.745 ;
      VIA 82.8 674.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 674.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 668.955 83.59 669.285 ;
      VIA 82.8 669.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 668.935 83.57 669.305 ;
      VIA 82.8 669.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 669.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 663.515 83.59 663.845 ;
      VIA 82.8 663.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 663.495 83.57 663.865 ;
      VIA 82.8 663.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 663.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 658.075 83.59 658.405 ;
      VIA 82.8 658.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 658.055 83.57 658.425 ;
      VIA 82.8 658.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 658.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 652.635 83.59 652.965 ;
      VIA 82.8 652.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 652.615 83.57 652.985 ;
      VIA 82.8 652.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 652.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 647.195 83.59 647.525 ;
      VIA 82.8 647.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 647.175 83.57 647.545 ;
      VIA 82.8 647.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 647.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 641.755 83.59 642.085 ;
      VIA 82.8 641.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 641.735 83.57 642.105 ;
      VIA 82.8 641.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 641.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 636.315 83.59 636.645 ;
      VIA 82.8 636.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 636.295 83.57 636.665 ;
      VIA 82.8 636.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 636.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 630.875 83.59 631.205 ;
      VIA 82.8 631.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 630.855 83.57 631.225 ;
      VIA 82.8 631.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 631.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 625.435 83.59 625.765 ;
      VIA 82.8 625.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 625.415 83.57 625.785 ;
      VIA 82.8 625.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 625.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 619.995 83.59 620.325 ;
      VIA 82.8 620.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 619.975 83.57 620.345 ;
      VIA 82.8 620.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 620.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 614.555 83.59 614.885 ;
      VIA 82.8 614.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 614.535 83.57 614.905 ;
      VIA 82.8 614.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 614.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 609.115 83.59 609.445 ;
      VIA 82.8 609.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 609.095 83.57 609.465 ;
      VIA 82.8 609.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 609.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 603.675 83.59 604.005 ;
      VIA 82.8 603.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 603.655 83.57 604.025 ;
      VIA 82.8 603.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 603.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 598.235 83.59 598.565 ;
      VIA 82.8 598.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 598.215 83.57 598.585 ;
      VIA 82.8 598.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 598.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 592.795 83.59 593.125 ;
      VIA 82.8 592.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 592.775 83.57 593.145 ;
      VIA 82.8 592.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 592.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 587.355 83.59 587.685 ;
      VIA 82.8 587.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 587.335 83.57 587.705 ;
      VIA 82.8 587.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 587.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 581.915 83.59 582.245 ;
      VIA 82.8 582.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 581.895 83.57 582.265 ;
      VIA 82.8 582.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 582.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 576.475 83.59 576.805 ;
      VIA 82.8 576.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 576.455 83.57 576.825 ;
      VIA 82.8 576.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 576.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 571.035 83.59 571.365 ;
      VIA 82.8 571.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 571.015 83.57 571.385 ;
      VIA 82.8 571.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 571.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 565.595 83.59 565.925 ;
      VIA 82.8 565.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 565.575 83.57 565.945 ;
      VIA 82.8 565.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 565.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 560.155 83.59 560.485 ;
      VIA 82.8 560.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 560.135 83.57 560.505 ;
      VIA 82.8 560.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 560.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 554.715 83.59 555.045 ;
      VIA 82.8 554.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 554.695 83.57 555.065 ;
      VIA 82.8 554.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 554.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 549.275 83.59 549.605 ;
      VIA 82.8 549.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 549.255 83.57 549.625 ;
      VIA 82.8 549.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 549.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 543.835 83.59 544.165 ;
      VIA 82.8 544 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 543.815 83.57 544.185 ;
      VIA 82.8 544 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 544 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 538.395 83.59 538.725 ;
      VIA 82.8 538.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 538.375 83.57 538.745 ;
      VIA 82.8 538.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 538.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 532.955 83.59 533.285 ;
      VIA 82.8 533.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 532.935 83.57 533.305 ;
      VIA 82.8 533.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 533.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 527.515 83.59 527.845 ;
      VIA 82.8 527.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 527.495 83.57 527.865 ;
      VIA 82.8 527.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 527.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 522.075 83.59 522.405 ;
      VIA 82.8 522.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 522.055 83.57 522.425 ;
      VIA 82.8 522.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 522.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 516.635 83.59 516.965 ;
      VIA 82.8 516.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 516.615 83.57 516.985 ;
      VIA 82.8 516.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 516.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 511.195 83.59 511.525 ;
      VIA 82.8 511.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 511.175 83.57 511.545 ;
      VIA 82.8 511.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 511.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 505.755 83.59 506.085 ;
      VIA 82.8 505.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 505.735 83.57 506.105 ;
      VIA 82.8 505.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 505.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 500.315 83.59 500.645 ;
      VIA 82.8 500.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 500.295 83.57 500.665 ;
      VIA 82.8 500.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 500.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 494.875 83.59 495.205 ;
      VIA 82.8 495.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 494.855 83.57 495.225 ;
      VIA 82.8 495.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 495.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 489.435 83.59 489.765 ;
      VIA 82.8 489.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 489.415 83.57 489.785 ;
      VIA 82.8 489.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 489.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 483.995 83.59 484.325 ;
      VIA 82.8 484.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 483.975 83.57 484.345 ;
      VIA 82.8 484.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 484.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 478.555 83.59 478.885 ;
      VIA 82.8 478.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 478.535 83.57 478.905 ;
      VIA 82.8 478.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 478.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 473.115 83.59 473.445 ;
      VIA 82.8 473.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 473.095 83.57 473.465 ;
      VIA 82.8 473.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 473.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 467.675 83.59 468.005 ;
      VIA 82.8 467.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 467.655 83.57 468.025 ;
      VIA 82.8 467.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 467.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 462.235 83.59 462.565 ;
      VIA 82.8 462.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 462.215 83.57 462.585 ;
      VIA 82.8 462.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 462.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 456.795 83.59 457.125 ;
      VIA 82.8 456.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 456.775 83.57 457.145 ;
      VIA 82.8 456.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 456.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 451.355 83.59 451.685 ;
      VIA 82.8 451.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 451.335 83.57 451.705 ;
      VIA 82.8 451.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 451.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 445.915 83.59 446.245 ;
      VIA 82.8 446.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 445.895 83.57 446.265 ;
      VIA 82.8 446.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 446.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 440.475 83.59 440.805 ;
      VIA 82.8 440.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 440.455 83.57 440.825 ;
      VIA 82.8 440.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 440.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 435.035 83.59 435.365 ;
      VIA 82.8 435.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 435.015 83.57 435.385 ;
      VIA 82.8 435.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 435.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 429.595 83.59 429.925 ;
      VIA 82.8 429.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 429.575 83.57 429.945 ;
      VIA 82.8 429.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 429.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 424.155 83.59 424.485 ;
      VIA 82.8 424.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 424.135 83.57 424.505 ;
      VIA 82.8 424.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 424.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 418.715 83.59 419.045 ;
      VIA 82.8 418.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 418.695 83.57 419.065 ;
      VIA 82.8 418.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 418.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 413.275 83.59 413.605 ;
      VIA 82.8 413.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 413.255 83.57 413.625 ;
      VIA 82.8 413.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 413.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 407.835 83.59 408.165 ;
      VIA 82.8 408 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 407.815 83.57 408.185 ;
      VIA 82.8 408 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 408 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 402.395 83.59 402.725 ;
      VIA 82.8 402.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 402.375 83.57 402.745 ;
      VIA 82.8 402.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 402.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 396.955 83.59 397.285 ;
      VIA 82.8 397.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 396.935 83.57 397.305 ;
      VIA 82.8 397.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 397.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 391.515 83.59 391.845 ;
      VIA 82.8 391.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 391.495 83.57 391.865 ;
      VIA 82.8 391.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 391.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 386.075 83.59 386.405 ;
      VIA 82.8 386.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 386.055 83.57 386.425 ;
      VIA 82.8 386.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 386.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 380.635 83.59 380.965 ;
      VIA 82.8 380.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 380.615 83.57 380.985 ;
      VIA 82.8 380.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 380.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 375.195 83.59 375.525 ;
      VIA 82.8 375.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 375.175 83.57 375.545 ;
      VIA 82.8 375.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 375.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 369.755 83.59 370.085 ;
      VIA 82.8 369.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 369.735 83.57 370.105 ;
      VIA 82.8 369.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 369.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 364.315 83.59 364.645 ;
      VIA 82.8 364.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 364.295 83.57 364.665 ;
      VIA 82.8 364.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 364.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 358.875 83.59 359.205 ;
      VIA 82.8 359.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 358.855 83.57 359.225 ;
      VIA 82.8 359.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 359.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 353.435 83.59 353.765 ;
      VIA 82.8 353.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 353.415 83.57 353.785 ;
      VIA 82.8 353.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 353.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 347.995 83.59 348.325 ;
      VIA 82.8 348.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 347.975 83.57 348.345 ;
      VIA 82.8 348.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 348.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 342.555 83.59 342.885 ;
      VIA 82.8 342.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 342.535 83.57 342.905 ;
      VIA 82.8 342.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 342.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 337.115 83.59 337.445 ;
      VIA 82.8 337.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 337.095 83.57 337.465 ;
      VIA 82.8 337.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 337.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 331.675 83.59 332.005 ;
      VIA 82.8 331.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 331.655 83.57 332.025 ;
      VIA 82.8 331.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 331.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 326.235 83.59 326.565 ;
      VIA 82.8 326.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 326.215 83.57 326.585 ;
      VIA 82.8 326.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 326.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 320.795 83.59 321.125 ;
      VIA 82.8 320.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 320.775 83.57 321.145 ;
      VIA 82.8 320.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 320.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 315.355 83.59 315.685 ;
      VIA 82.8 315.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 315.335 83.57 315.705 ;
      VIA 82.8 315.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 315.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 309.915 83.59 310.245 ;
      VIA 82.8 310.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 309.895 83.57 310.265 ;
      VIA 82.8 310.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 310.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 304.475 83.59 304.805 ;
      VIA 82.8 304.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 304.455 83.57 304.825 ;
      VIA 82.8 304.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 304.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 299.035 83.59 299.365 ;
      VIA 82.8 299.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 299.015 83.57 299.385 ;
      VIA 82.8 299.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 299.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 293.595 83.59 293.925 ;
      VIA 82.8 293.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 293.575 83.57 293.945 ;
      VIA 82.8 293.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 293.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 288.155 83.59 288.485 ;
      VIA 82.8 288.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 288.135 83.57 288.505 ;
      VIA 82.8 288.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 288.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 282.715 83.59 283.045 ;
      VIA 82.8 282.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 282.695 83.57 283.065 ;
      VIA 82.8 282.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 282.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 277.275 83.59 277.605 ;
      VIA 82.8 277.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 277.255 83.57 277.625 ;
      VIA 82.8 277.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 277.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 271.835 83.59 272.165 ;
      VIA 82.8 272 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 271.815 83.57 272.185 ;
      VIA 82.8 272 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 272 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 266.395 83.59 266.725 ;
      VIA 82.8 266.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 266.375 83.57 266.745 ;
      VIA 82.8 266.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 266.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 260.955 83.59 261.285 ;
      VIA 82.8 261.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 260.935 83.57 261.305 ;
      VIA 82.8 261.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 261.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 255.515 83.59 255.845 ;
      VIA 82.8 255.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 255.495 83.57 255.865 ;
      VIA 82.8 255.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 255.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 250.075 83.59 250.405 ;
      VIA 82.8 250.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 250.055 83.57 250.425 ;
      VIA 82.8 250.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 250.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 244.635 83.59 244.965 ;
      VIA 82.8 244.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 244.615 83.57 244.985 ;
      VIA 82.8 244.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 244.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 239.195 83.59 239.525 ;
      VIA 82.8 239.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 239.175 83.57 239.545 ;
      VIA 82.8 239.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 239.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 233.755 83.59 234.085 ;
      VIA 82.8 233.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 233.735 83.57 234.105 ;
      VIA 82.8 233.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 233.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 228.315 83.59 228.645 ;
      VIA 82.8 228.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 228.295 83.57 228.665 ;
      VIA 82.8 228.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 228.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 222.875 83.59 223.205 ;
      VIA 82.8 223.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 222.855 83.57 223.225 ;
      VIA 82.8 223.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 223.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 217.435 83.59 217.765 ;
      VIA 82.8 217.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 217.415 83.57 217.785 ;
      VIA 82.8 217.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 217.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 211.995 83.59 212.325 ;
      VIA 82.8 212.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 211.975 83.57 212.345 ;
      VIA 82.8 212.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 212.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 206.555 83.59 206.885 ;
      VIA 82.8 206.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 206.535 83.57 206.905 ;
      VIA 82.8 206.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 206.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 201.115 83.59 201.445 ;
      VIA 82.8 201.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 201.095 83.57 201.465 ;
      VIA 82.8 201.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 201.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 195.675 83.59 196.005 ;
      VIA 82.8 195.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 195.655 83.57 196.025 ;
      VIA 82.8 195.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 195.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 190.235 83.59 190.565 ;
      VIA 82.8 190.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 190.215 83.57 190.585 ;
      VIA 82.8 190.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 190.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 184.795 83.59 185.125 ;
      VIA 82.8 184.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 184.775 83.57 185.145 ;
      VIA 82.8 184.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 184.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 179.355 83.59 179.685 ;
      VIA 82.8 179.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 179.335 83.57 179.705 ;
      VIA 82.8 179.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 179.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 173.915 83.59 174.245 ;
      VIA 82.8 174.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 173.895 83.57 174.265 ;
      VIA 82.8 174.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 174.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 168.475 83.59 168.805 ;
      VIA 82.8 168.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 168.455 83.57 168.825 ;
      VIA 82.8 168.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 168.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 163.035 83.59 163.365 ;
      VIA 82.8 163.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 163.015 83.57 163.385 ;
      VIA 82.8 163.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 163.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 157.595 83.59 157.925 ;
      VIA 82.8 157.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 157.575 83.57 157.945 ;
      VIA 82.8 157.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 157.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 152.155 83.59 152.485 ;
      VIA 82.8 152.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 152.135 83.57 152.505 ;
      VIA 82.8 152.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 152.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 146.715 83.59 147.045 ;
      VIA 82.8 146.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 146.695 83.57 147.065 ;
      VIA 82.8 146.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 146.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 141.275 83.59 141.605 ;
      VIA 82.8 141.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 141.255 83.57 141.625 ;
      VIA 82.8 141.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 141.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 135.835 83.59 136.165 ;
      VIA 82.8 136 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 135.815 83.57 136.185 ;
      VIA 82.8 136 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 136 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 130.395 83.59 130.725 ;
      VIA 82.8 130.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 130.375 83.57 130.745 ;
      VIA 82.8 130.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 130.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 124.955 83.59 125.285 ;
      VIA 82.8 125.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 124.935 83.57 125.305 ;
      VIA 82.8 125.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 125.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 119.515 83.59 119.845 ;
      VIA 82.8 119.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 119.495 83.57 119.865 ;
      VIA 82.8 119.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 119.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 114.075 83.59 114.405 ;
      VIA 82.8 114.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 114.055 83.57 114.425 ;
      VIA 82.8 114.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 114.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 108.635 83.59 108.965 ;
      VIA 82.8 108.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 108.615 83.57 108.985 ;
      VIA 82.8 108.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 108.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 103.195 83.59 103.525 ;
      VIA 82.8 103.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 103.175 83.57 103.545 ;
      VIA 82.8 103.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 103.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 97.755 83.59 98.085 ;
      VIA 82.8 97.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 97.735 83.57 98.105 ;
      VIA 82.8 97.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 97.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 92.315 83.59 92.645 ;
      VIA 82.8 92.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 92.295 83.57 92.665 ;
      VIA 82.8 92.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 92.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 86.875 83.59 87.205 ;
      VIA 82.8 87.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 86.855 83.57 87.225 ;
      VIA 82.8 87.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 87.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 81.435 83.59 81.765 ;
      VIA 82.8 81.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 81.415 83.57 81.785 ;
      VIA 82.8 81.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 81.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 75.995 83.59 76.325 ;
      VIA 82.8 76.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 75.975 83.57 76.345 ;
      VIA 82.8 76.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 76.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 70.555 83.59 70.885 ;
      VIA 82.8 70.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 70.535 83.57 70.905 ;
      VIA 82.8 70.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 70.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 65.115 83.59 65.445 ;
      VIA 82.8 65.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 65.095 83.57 65.465 ;
      VIA 82.8 65.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 65.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 59.675 83.59 60.005 ;
      VIA 82.8 59.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 59.655 83.57 60.025 ;
      VIA 82.8 59.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 59.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 54.235 83.59 54.565 ;
      VIA 82.8 54.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 54.215 83.57 54.585 ;
      VIA 82.8 54.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 54.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 48.795 83.59 49.125 ;
      VIA 82.8 48.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 48.775 83.57 49.145 ;
      VIA 82.8 48.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 48.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 43.355 83.59 43.685 ;
      VIA 82.8 43.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 43.335 83.57 43.705 ;
      VIA 82.8 43.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 43.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 37.915 83.59 38.245 ;
      VIA 82.8 38.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 37.895 83.57 38.265 ;
      VIA 82.8 38.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 38.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 32.475 83.59 32.805 ;
      VIA 82.8 32.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 32.455 83.57 32.825 ;
      VIA 82.8 32.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 32.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 27.035 83.59 27.365 ;
      VIA 82.8 27.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 27.015 83.57 27.385 ;
      VIA 82.8 27.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 27.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 21.595 83.59 21.925 ;
      VIA 82.8 21.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 21.575 83.57 21.945 ;
      VIA 82.8 21.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 21.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 16.155 83.59 16.485 ;
      VIA 82.8 16.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 16.135 83.57 16.505 ;
      VIA 82.8 16.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 16.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 10.715 83.59 11.045 ;
      VIA 82.8 10.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 10.695 83.57 11.065 ;
      VIA 82.8 10.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 10.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  82.01 5.275 83.59 5.605 ;
      VIA 82.8 5.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  82.03 5.255 83.57 5.625 ;
      VIA 82.8 5.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 82.8 5.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 701.595 56.45 701.925 ;
      VIA 55.66 701.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 701.575 56.43 701.945 ;
      VIA 55.66 701.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 701.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 696.155 56.45 696.485 ;
      VIA 55.66 696.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 696.135 56.43 696.505 ;
      VIA 55.66 696.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 696.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 690.715 56.45 691.045 ;
      VIA 55.66 690.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 690.695 56.43 691.065 ;
      VIA 55.66 690.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 690.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 685.275 56.45 685.605 ;
      VIA 55.66 685.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 685.255 56.43 685.625 ;
      VIA 55.66 685.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 685.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 679.835 56.45 680.165 ;
      VIA 55.66 680 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 679.815 56.43 680.185 ;
      VIA 55.66 680 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 680 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 674.395 56.45 674.725 ;
      VIA 55.66 674.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 674.375 56.43 674.745 ;
      VIA 55.66 674.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 674.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 668.955 56.45 669.285 ;
      VIA 55.66 669.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 668.935 56.43 669.305 ;
      VIA 55.66 669.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 669.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 663.515 56.45 663.845 ;
      VIA 55.66 663.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 663.495 56.43 663.865 ;
      VIA 55.66 663.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 663.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 658.075 56.45 658.405 ;
      VIA 55.66 658.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 658.055 56.43 658.425 ;
      VIA 55.66 658.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 658.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 652.635 56.45 652.965 ;
      VIA 55.66 652.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 652.615 56.43 652.985 ;
      VIA 55.66 652.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 652.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 647.195 56.45 647.525 ;
      VIA 55.66 647.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 647.175 56.43 647.545 ;
      VIA 55.66 647.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 647.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 641.755 56.45 642.085 ;
      VIA 55.66 641.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 641.735 56.43 642.105 ;
      VIA 55.66 641.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 641.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 636.315 56.45 636.645 ;
      VIA 55.66 636.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 636.295 56.43 636.665 ;
      VIA 55.66 636.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 636.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 630.875 56.45 631.205 ;
      VIA 55.66 631.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 630.855 56.43 631.225 ;
      VIA 55.66 631.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 631.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 625.435 56.45 625.765 ;
      VIA 55.66 625.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 625.415 56.43 625.785 ;
      VIA 55.66 625.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 625.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 619.995 56.45 620.325 ;
      VIA 55.66 620.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 619.975 56.43 620.345 ;
      VIA 55.66 620.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 620.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 614.555 56.45 614.885 ;
      VIA 55.66 614.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 614.535 56.43 614.905 ;
      VIA 55.66 614.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 614.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 609.115 56.45 609.445 ;
      VIA 55.66 609.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 609.095 56.43 609.465 ;
      VIA 55.66 609.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 609.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 603.675 56.45 604.005 ;
      VIA 55.66 603.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 603.655 56.43 604.025 ;
      VIA 55.66 603.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 603.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 598.235 56.45 598.565 ;
      VIA 55.66 598.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 598.215 56.43 598.585 ;
      VIA 55.66 598.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 598.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 592.795 56.45 593.125 ;
      VIA 55.66 592.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 592.775 56.43 593.145 ;
      VIA 55.66 592.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 592.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 587.355 56.45 587.685 ;
      VIA 55.66 587.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 587.335 56.43 587.705 ;
      VIA 55.66 587.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 587.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 581.915 56.45 582.245 ;
      VIA 55.66 582.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 581.895 56.43 582.265 ;
      VIA 55.66 582.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 582.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 576.475 56.45 576.805 ;
      VIA 55.66 576.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 576.455 56.43 576.825 ;
      VIA 55.66 576.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 576.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 571.035 56.45 571.365 ;
      VIA 55.66 571.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 571.015 56.43 571.385 ;
      VIA 55.66 571.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 571.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 565.595 56.45 565.925 ;
      VIA 55.66 565.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 565.575 56.43 565.945 ;
      VIA 55.66 565.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 565.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 560.155 56.45 560.485 ;
      VIA 55.66 560.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 560.135 56.43 560.505 ;
      VIA 55.66 560.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 560.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 554.715 56.45 555.045 ;
      VIA 55.66 554.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 554.695 56.43 555.065 ;
      VIA 55.66 554.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 554.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 549.275 56.45 549.605 ;
      VIA 55.66 549.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 549.255 56.43 549.625 ;
      VIA 55.66 549.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 549.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 543.835 56.45 544.165 ;
      VIA 55.66 544 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 543.815 56.43 544.185 ;
      VIA 55.66 544 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 544 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 538.395 56.45 538.725 ;
      VIA 55.66 538.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 538.375 56.43 538.745 ;
      VIA 55.66 538.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 538.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 532.955 56.45 533.285 ;
      VIA 55.66 533.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 532.935 56.43 533.305 ;
      VIA 55.66 533.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 533.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 527.515 56.45 527.845 ;
      VIA 55.66 527.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 527.495 56.43 527.865 ;
      VIA 55.66 527.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 527.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 522.075 56.45 522.405 ;
      VIA 55.66 522.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 522.055 56.43 522.425 ;
      VIA 55.66 522.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 522.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 516.635 56.45 516.965 ;
      VIA 55.66 516.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 516.615 56.43 516.985 ;
      VIA 55.66 516.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 516.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 511.195 56.45 511.525 ;
      VIA 55.66 511.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 511.175 56.43 511.545 ;
      VIA 55.66 511.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 511.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 505.755 56.45 506.085 ;
      VIA 55.66 505.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 505.735 56.43 506.105 ;
      VIA 55.66 505.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 505.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 500.315 56.45 500.645 ;
      VIA 55.66 500.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 500.295 56.43 500.665 ;
      VIA 55.66 500.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 500.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 494.875 56.45 495.205 ;
      VIA 55.66 495.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 494.855 56.43 495.225 ;
      VIA 55.66 495.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 495.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 489.435 56.45 489.765 ;
      VIA 55.66 489.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 489.415 56.43 489.785 ;
      VIA 55.66 489.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 489.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 483.995 56.45 484.325 ;
      VIA 55.66 484.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 483.975 56.43 484.345 ;
      VIA 55.66 484.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 484.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 478.555 56.45 478.885 ;
      VIA 55.66 478.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 478.535 56.43 478.905 ;
      VIA 55.66 478.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 478.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 473.115 56.45 473.445 ;
      VIA 55.66 473.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 473.095 56.43 473.465 ;
      VIA 55.66 473.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 473.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 467.675 56.45 468.005 ;
      VIA 55.66 467.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 467.655 56.43 468.025 ;
      VIA 55.66 467.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 467.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 462.235 56.45 462.565 ;
      VIA 55.66 462.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 462.215 56.43 462.585 ;
      VIA 55.66 462.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 462.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 456.795 56.45 457.125 ;
      VIA 55.66 456.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 456.775 56.43 457.145 ;
      VIA 55.66 456.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 456.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 451.355 56.45 451.685 ;
      VIA 55.66 451.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 451.335 56.43 451.705 ;
      VIA 55.66 451.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 451.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 445.915 56.45 446.245 ;
      VIA 55.66 446.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 445.895 56.43 446.265 ;
      VIA 55.66 446.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 446.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 440.475 56.45 440.805 ;
      VIA 55.66 440.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 440.455 56.43 440.825 ;
      VIA 55.66 440.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 440.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 435.035 56.45 435.365 ;
      VIA 55.66 435.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 435.015 56.43 435.385 ;
      VIA 55.66 435.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 435.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 429.595 56.45 429.925 ;
      VIA 55.66 429.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 429.575 56.43 429.945 ;
      VIA 55.66 429.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 429.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 424.155 56.45 424.485 ;
      VIA 55.66 424.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 424.135 56.43 424.505 ;
      VIA 55.66 424.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 424.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 418.715 56.45 419.045 ;
      VIA 55.66 418.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 418.695 56.43 419.065 ;
      VIA 55.66 418.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 418.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 413.275 56.45 413.605 ;
      VIA 55.66 413.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 413.255 56.43 413.625 ;
      VIA 55.66 413.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 413.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 407.835 56.45 408.165 ;
      VIA 55.66 408 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 407.815 56.43 408.185 ;
      VIA 55.66 408 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 408 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 402.395 56.45 402.725 ;
      VIA 55.66 402.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 402.375 56.43 402.745 ;
      VIA 55.66 402.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 402.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 396.955 56.45 397.285 ;
      VIA 55.66 397.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 396.935 56.43 397.305 ;
      VIA 55.66 397.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 397.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 391.515 56.45 391.845 ;
      VIA 55.66 391.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 391.495 56.43 391.865 ;
      VIA 55.66 391.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 391.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 386.075 56.45 386.405 ;
      VIA 55.66 386.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 386.055 56.43 386.425 ;
      VIA 55.66 386.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 386.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 380.635 56.45 380.965 ;
      VIA 55.66 380.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 380.615 56.43 380.985 ;
      VIA 55.66 380.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 380.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 375.195 56.45 375.525 ;
      VIA 55.66 375.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 375.175 56.43 375.545 ;
      VIA 55.66 375.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 375.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 369.755 56.45 370.085 ;
      VIA 55.66 369.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 369.735 56.43 370.105 ;
      VIA 55.66 369.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 369.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 364.315 56.45 364.645 ;
      VIA 55.66 364.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 364.295 56.43 364.665 ;
      VIA 55.66 364.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 364.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 358.875 56.45 359.205 ;
      VIA 55.66 359.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 358.855 56.43 359.225 ;
      VIA 55.66 359.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 359.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 353.435 56.45 353.765 ;
      VIA 55.66 353.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 353.415 56.43 353.785 ;
      VIA 55.66 353.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 353.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 347.995 56.45 348.325 ;
      VIA 55.66 348.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 347.975 56.43 348.345 ;
      VIA 55.66 348.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 348.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 342.555 56.45 342.885 ;
      VIA 55.66 342.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 342.535 56.43 342.905 ;
      VIA 55.66 342.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 342.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 337.115 56.45 337.445 ;
      VIA 55.66 337.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 337.095 56.43 337.465 ;
      VIA 55.66 337.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 337.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 331.675 56.45 332.005 ;
      VIA 55.66 331.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 331.655 56.43 332.025 ;
      VIA 55.66 331.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 331.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 326.235 56.45 326.565 ;
      VIA 55.66 326.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 326.215 56.43 326.585 ;
      VIA 55.66 326.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 326.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 320.795 56.45 321.125 ;
      VIA 55.66 320.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 320.775 56.43 321.145 ;
      VIA 55.66 320.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 320.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 315.355 56.45 315.685 ;
      VIA 55.66 315.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 315.335 56.43 315.705 ;
      VIA 55.66 315.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 315.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 309.915 56.45 310.245 ;
      VIA 55.66 310.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 309.895 56.43 310.265 ;
      VIA 55.66 310.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 310.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 304.475 56.45 304.805 ;
      VIA 55.66 304.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 304.455 56.43 304.825 ;
      VIA 55.66 304.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 304.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 299.035 56.45 299.365 ;
      VIA 55.66 299.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 299.015 56.43 299.385 ;
      VIA 55.66 299.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 299.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 293.595 56.45 293.925 ;
      VIA 55.66 293.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 293.575 56.43 293.945 ;
      VIA 55.66 293.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 293.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 288.155 56.45 288.485 ;
      VIA 55.66 288.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 288.135 56.43 288.505 ;
      VIA 55.66 288.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 288.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 282.715 56.45 283.045 ;
      VIA 55.66 282.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 282.695 56.43 283.065 ;
      VIA 55.66 282.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 282.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 277.275 56.45 277.605 ;
      VIA 55.66 277.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 277.255 56.43 277.625 ;
      VIA 55.66 277.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 277.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 271.835 56.45 272.165 ;
      VIA 55.66 272 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 271.815 56.43 272.185 ;
      VIA 55.66 272 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 272 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 266.395 56.45 266.725 ;
      VIA 55.66 266.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 266.375 56.43 266.745 ;
      VIA 55.66 266.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 266.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 260.955 56.45 261.285 ;
      VIA 55.66 261.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 260.935 56.43 261.305 ;
      VIA 55.66 261.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 261.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 255.515 56.45 255.845 ;
      VIA 55.66 255.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 255.495 56.43 255.865 ;
      VIA 55.66 255.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 255.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 250.075 56.45 250.405 ;
      VIA 55.66 250.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 250.055 56.43 250.425 ;
      VIA 55.66 250.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 250.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 244.635 56.45 244.965 ;
      VIA 55.66 244.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 244.615 56.43 244.985 ;
      VIA 55.66 244.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 244.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 239.195 56.45 239.525 ;
      VIA 55.66 239.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 239.175 56.43 239.545 ;
      VIA 55.66 239.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 239.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 233.755 56.45 234.085 ;
      VIA 55.66 233.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 233.735 56.43 234.105 ;
      VIA 55.66 233.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 233.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 228.315 56.45 228.645 ;
      VIA 55.66 228.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 228.295 56.43 228.665 ;
      VIA 55.66 228.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 228.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 222.875 56.45 223.205 ;
      VIA 55.66 223.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 222.855 56.43 223.225 ;
      VIA 55.66 223.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 223.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 217.435 56.45 217.765 ;
      VIA 55.66 217.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 217.415 56.43 217.785 ;
      VIA 55.66 217.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 217.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 211.995 56.45 212.325 ;
      VIA 55.66 212.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 211.975 56.43 212.345 ;
      VIA 55.66 212.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 212.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 206.555 56.45 206.885 ;
      VIA 55.66 206.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 206.535 56.43 206.905 ;
      VIA 55.66 206.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 206.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 201.115 56.45 201.445 ;
      VIA 55.66 201.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 201.095 56.43 201.465 ;
      VIA 55.66 201.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 201.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 195.675 56.45 196.005 ;
      VIA 55.66 195.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 195.655 56.43 196.025 ;
      VIA 55.66 195.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 195.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 190.235 56.45 190.565 ;
      VIA 55.66 190.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 190.215 56.43 190.585 ;
      VIA 55.66 190.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 190.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 184.795 56.45 185.125 ;
      VIA 55.66 184.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 184.775 56.43 185.145 ;
      VIA 55.66 184.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 184.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 179.355 56.45 179.685 ;
      VIA 55.66 179.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 179.335 56.43 179.705 ;
      VIA 55.66 179.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 179.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 173.915 56.45 174.245 ;
      VIA 55.66 174.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 173.895 56.43 174.265 ;
      VIA 55.66 174.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 174.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 168.475 56.45 168.805 ;
      VIA 55.66 168.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 168.455 56.43 168.825 ;
      VIA 55.66 168.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 168.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 163.035 56.45 163.365 ;
      VIA 55.66 163.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 163.015 56.43 163.385 ;
      VIA 55.66 163.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 163.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 157.595 56.45 157.925 ;
      VIA 55.66 157.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 157.575 56.43 157.945 ;
      VIA 55.66 157.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 157.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 152.155 56.45 152.485 ;
      VIA 55.66 152.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 152.135 56.43 152.505 ;
      VIA 55.66 152.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 152.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 146.715 56.45 147.045 ;
      VIA 55.66 146.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 146.695 56.43 147.065 ;
      VIA 55.66 146.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 146.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 141.275 56.45 141.605 ;
      VIA 55.66 141.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 141.255 56.43 141.625 ;
      VIA 55.66 141.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 141.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 135.835 56.45 136.165 ;
      VIA 55.66 136 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 135.815 56.43 136.185 ;
      VIA 55.66 136 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 136 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 130.395 56.45 130.725 ;
      VIA 55.66 130.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 130.375 56.43 130.745 ;
      VIA 55.66 130.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 130.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 124.955 56.45 125.285 ;
      VIA 55.66 125.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 124.935 56.43 125.305 ;
      VIA 55.66 125.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 125.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 119.515 56.45 119.845 ;
      VIA 55.66 119.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 119.495 56.43 119.865 ;
      VIA 55.66 119.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 119.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 114.075 56.45 114.405 ;
      VIA 55.66 114.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 114.055 56.43 114.425 ;
      VIA 55.66 114.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 114.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 108.635 56.45 108.965 ;
      VIA 55.66 108.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 108.615 56.43 108.985 ;
      VIA 55.66 108.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 108.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 103.195 56.45 103.525 ;
      VIA 55.66 103.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 103.175 56.43 103.545 ;
      VIA 55.66 103.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 103.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 97.755 56.45 98.085 ;
      VIA 55.66 97.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 97.735 56.43 98.105 ;
      VIA 55.66 97.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 97.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 92.315 56.45 92.645 ;
      VIA 55.66 92.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 92.295 56.43 92.665 ;
      VIA 55.66 92.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 92.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 86.875 56.45 87.205 ;
      VIA 55.66 87.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 86.855 56.43 87.225 ;
      VIA 55.66 87.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 87.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 81.435 56.45 81.765 ;
      VIA 55.66 81.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 81.415 56.43 81.785 ;
      VIA 55.66 81.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 81.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 75.995 56.45 76.325 ;
      VIA 55.66 76.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 75.975 56.43 76.345 ;
      VIA 55.66 76.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 76.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 70.555 56.45 70.885 ;
      VIA 55.66 70.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 70.535 56.43 70.905 ;
      VIA 55.66 70.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 70.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 65.115 56.45 65.445 ;
      VIA 55.66 65.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 65.095 56.43 65.465 ;
      VIA 55.66 65.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 65.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 59.675 56.45 60.005 ;
      VIA 55.66 59.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 59.655 56.43 60.025 ;
      VIA 55.66 59.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 59.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 54.235 56.45 54.565 ;
      VIA 55.66 54.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 54.215 56.43 54.585 ;
      VIA 55.66 54.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 54.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 48.795 56.45 49.125 ;
      VIA 55.66 48.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 48.775 56.43 49.145 ;
      VIA 55.66 48.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 48.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 43.355 56.45 43.685 ;
      VIA 55.66 43.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 43.335 56.43 43.705 ;
      VIA 55.66 43.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 43.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 37.915 56.45 38.245 ;
      VIA 55.66 38.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 37.895 56.43 38.265 ;
      VIA 55.66 38.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 38.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 32.475 56.45 32.805 ;
      VIA 55.66 32.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 32.455 56.43 32.825 ;
      VIA 55.66 32.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 32.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 27.035 56.45 27.365 ;
      VIA 55.66 27.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 27.015 56.43 27.385 ;
      VIA 55.66 27.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 27.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 21.595 56.45 21.925 ;
      VIA 55.66 21.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 21.575 56.43 21.945 ;
      VIA 55.66 21.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 21.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 16.155 56.45 16.485 ;
      VIA 55.66 16.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 16.135 56.43 16.505 ;
      VIA 55.66 16.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 16.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 10.715 56.45 11.045 ;
      VIA 55.66 10.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 10.695 56.43 11.065 ;
      VIA 55.66 10.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 10.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  54.87 5.275 56.45 5.605 ;
      VIA 55.66 5.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  54.89 5.255 56.43 5.625 ;
      VIA 55.66 5.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 55.66 5.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 701.595 29.31 701.925 ;
      VIA 28.52 701.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 701.575 29.29 701.945 ;
      VIA 28.52 701.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 701.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 696.155 29.31 696.485 ;
      VIA 28.52 696.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 696.135 29.29 696.505 ;
      VIA 28.52 696.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 696.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 690.715 29.31 691.045 ;
      VIA 28.52 690.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 690.695 29.29 691.065 ;
      VIA 28.52 690.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 690.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 685.275 29.31 685.605 ;
      VIA 28.52 685.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 685.255 29.29 685.625 ;
      VIA 28.52 685.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 685.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 679.835 29.31 680.165 ;
      VIA 28.52 680 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 679.815 29.29 680.185 ;
      VIA 28.52 680 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 680 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 674.395 29.31 674.725 ;
      VIA 28.52 674.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 674.375 29.29 674.745 ;
      VIA 28.52 674.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 674.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 668.955 29.31 669.285 ;
      VIA 28.52 669.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 668.935 29.29 669.305 ;
      VIA 28.52 669.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 669.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 663.515 29.31 663.845 ;
      VIA 28.52 663.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 663.495 29.29 663.865 ;
      VIA 28.52 663.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 663.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 658.075 29.31 658.405 ;
      VIA 28.52 658.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 658.055 29.29 658.425 ;
      VIA 28.52 658.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 658.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 652.635 29.31 652.965 ;
      VIA 28.52 652.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 652.615 29.29 652.985 ;
      VIA 28.52 652.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 652.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 647.195 29.31 647.525 ;
      VIA 28.52 647.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 647.175 29.29 647.545 ;
      VIA 28.52 647.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 647.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 641.755 29.31 642.085 ;
      VIA 28.52 641.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 641.735 29.29 642.105 ;
      VIA 28.52 641.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 641.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 636.315 29.31 636.645 ;
      VIA 28.52 636.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 636.295 29.29 636.665 ;
      VIA 28.52 636.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 636.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 630.875 29.31 631.205 ;
      VIA 28.52 631.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 630.855 29.29 631.225 ;
      VIA 28.52 631.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 631.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 625.435 29.31 625.765 ;
      VIA 28.52 625.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 625.415 29.29 625.785 ;
      VIA 28.52 625.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 625.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 619.995 29.31 620.325 ;
      VIA 28.52 620.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 619.975 29.29 620.345 ;
      VIA 28.52 620.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 620.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 614.555 29.31 614.885 ;
      VIA 28.52 614.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 614.535 29.29 614.905 ;
      VIA 28.52 614.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 614.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 609.115 29.31 609.445 ;
      VIA 28.52 609.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 609.095 29.29 609.465 ;
      VIA 28.52 609.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 609.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 603.675 29.31 604.005 ;
      VIA 28.52 603.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 603.655 29.29 604.025 ;
      VIA 28.52 603.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 603.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 598.235 29.31 598.565 ;
      VIA 28.52 598.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 598.215 29.29 598.585 ;
      VIA 28.52 598.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 598.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 592.795 29.31 593.125 ;
      VIA 28.52 592.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 592.775 29.29 593.145 ;
      VIA 28.52 592.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 592.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 587.355 29.31 587.685 ;
      VIA 28.52 587.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 587.335 29.29 587.705 ;
      VIA 28.52 587.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 587.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 581.915 29.31 582.245 ;
      VIA 28.52 582.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 581.895 29.29 582.265 ;
      VIA 28.52 582.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 582.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 576.475 29.31 576.805 ;
      VIA 28.52 576.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 576.455 29.29 576.825 ;
      VIA 28.52 576.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 576.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 571.035 29.31 571.365 ;
      VIA 28.52 571.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 571.015 29.29 571.385 ;
      VIA 28.52 571.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 571.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 565.595 29.31 565.925 ;
      VIA 28.52 565.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 565.575 29.29 565.945 ;
      VIA 28.52 565.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 565.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 560.155 29.31 560.485 ;
      VIA 28.52 560.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 560.135 29.29 560.505 ;
      VIA 28.52 560.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 560.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 554.715 29.31 555.045 ;
      VIA 28.52 554.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 554.695 29.29 555.065 ;
      VIA 28.52 554.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 554.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 549.275 29.31 549.605 ;
      VIA 28.52 549.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 549.255 29.29 549.625 ;
      VIA 28.52 549.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 549.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 543.835 29.31 544.165 ;
      VIA 28.52 544 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 543.815 29.29 544.185 ;
      VIA 28.52 544 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 544 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 538.395 29.31 538.725 ;
      VIA 28.52 538.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 538.375 29.29 538.745 ;
      VIA 28.52 538.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 538.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 532.955 29.31 533.285 ;
      VIA 28.52 533.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 532.935 29.29 533.305 ;
      VIA 28.52 533.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 533.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 527.515 29.31 527.845 ;
      VIA 28.52 527.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 527.495 29.29 527.865 ;
      VIA 28.52 527.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 527.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 522.075 29.31 522.405 ;
      VIA 28.52 522.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 522.055 29.29 522.425 ;
      VIA 28.52 522.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 522.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 516.635 29.31 516.965 ;
      VIA 28.52 516.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 516.615 29.29 516.985 ;
      VIA 28.52 516.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 516.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 511.195 29.31 511.525 ;
      VIA 28.52 511.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 511.175 29.29 511.545 ;
      VIA 28.52 511.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 511.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 505.755 29.31 506.085 ;
      VIA 28.52 505.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 505.735 29.29 506.105 ;
      VIA 28.52 505.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 505.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 500.315 29.31 500.645 ;
      VIA 28.52 500.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 500.295 29.29 500.665 ;
      VIA 28.52 500.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 500.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 494.875 29.31 495.205 ;
      VIA 28.52 495.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 494.855 29.29 495.225 ;
      VIA 28.52 495.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 495.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 489.435 29.31 489.765 ;
      VIA 28.52 489.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 489.415 29.29 489.785 ;
      VIA 28.52 489.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 489.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 483.995 29.31 484.325 ;
      VIA 28.52 484.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 483.975 29.29 484.345 ;
      VIA 28.52 484.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 484.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 478.555 29.31 478.885 ;
      VIA 28.52 478.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 478.535 29.29 478.905 ;
      VIA 28.52 478.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 478.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 473.115 29.31 473.445 ;
      VIA 28.52 473.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 473.095 29.29 473.465 ;
      VIA 28.52 473.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 473.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 467.675 29.31 468.005 ;
      VIA 28.52 467.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 467.655 29.29 468.025 ;
      VIA 28.52 467.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 467.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 462.235 29.31 462.565 ;
      VIA 28.52 462.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 462.215 29.29 462.585 ;
      VIA 28.52 462.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 462.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 456.795 29.31 457.125 ;
      VIA 28.52 456.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 456.775 29.29 457.145 ;
      VIA 28.52 456.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 456.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 451.355 29.31 451.685 ;
      VIA 28.52 451.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 451.335 29.29 451.705 ;
      VIA 28.52 451.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 451.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 445.915 29.31 446.245 ;
      VIA 28.52 446.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 445.895 29.29 446.265 ;
      VIA 28.52 446.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 446.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 440.475 29.31 440.805 ;
      VIA 28.52 440.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 440.455 29.29 440.825 ;
      VIA 28.52 440.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 440.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 435.035 29.31 435.365 ;
      VIA 28.52 435.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 435.015 29.29 435.385 ;
      VIA 28.52 435.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 435.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 429.595 29.31 429.925 ;
      VIA 28.52 429.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 429.575 29.29 429.945 ;
      VIA 28.52 429.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 429.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 424.155 29.31 424.485 ;
      VIA 28.52 424.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 424.135 29.29 424.505 ;
      VIA 28.52 424.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 424.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 418.715 29.31 419.045 ;
      VIA 28.52 418.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 418.695 29.29 419.065 ;
      VIA 28.52 418.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 418.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 413.275 29.31 413.605 ;
      VIA 28.52 413.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 413.255 29.29 413.625 ;
      VIA 28.52 413.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 413.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 407.835 29.31 408.165 ;
      VIA 28.52 408 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 407.815 29.29 408.185 ;
      VIA 28.52 408 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 408 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 402.395 29.31 402.725 ;
      VIA 28.52 402.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 402.375 29.29 402.745 ;
      VIA 28.52 402.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 402.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 396.955 29.31 397.285 ;
      VIA 28.52 397.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 396.935 29.29 397.305 ;
      VIA 28.52 397.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 397.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 391.515 29.31 391.845 ;
      VIA 28.52 391.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 391.495 29.29 391.865 ;
      VIA 28.52 391.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 391.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 386.075 29.31 386.405 ;
      VIA 28.52 386.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 386.055 29.29 386.425 ;
      VIA 28.52 386.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 386.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 380.635 29.31 380.965 ;
      VIA 28.52 380.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 380.615 29.29 380.985 ;
      VIA 28.52 380.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 380.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 375.195 29.31 375.525 ;
      VIA 28.52 375.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 375.175 29.29 375.545 ;
      VIA 28.52 375.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 375.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 369.755 29.31 370.085 ;
      VIA 28.52 369.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 369.735 29.29 370.105 ;
      VIA 28.52 369.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 369.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 364.315 29.31 364.645 ;
      VIA 28.52 364.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 364.295 29.29 364.665 ;
      VIA 28.52 364.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 364.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 358.875 29.31 359.205 ;
      VIA 28.52 359.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 358.855 29.29 359.225 ;
      VIA 28.52 359.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 359.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 353.435 29.31 353.765 ;
      VIA 28.52 353.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 353.415 29.29 353.785 ;
      VIA 28.52 353.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 353.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 347.995 29.31 348.325 ;
      VIA 28.52 348.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 347.975 29.29 348.345 ;
      VIA 28.52 348.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 348.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 342.555 29.31 342.885 ;
      VIA 28.52 342.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 342.535 29.29 342.905 ;
      VIA 28.52 342.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 342.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 337.115 29.31 337.445 ;
      VIA 28.52 337.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 337.095 29.29 337.465 ;
      VIA 28.52 337.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 337.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 331.675 29.31 332.005 ;
      VIA 28.52 331.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 331.655 29.29 332.025 ;
      VIA 28.52 331.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 331.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 326.235 29.31 326.565 ;
      VIA 28.52 326.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 326.215 29.29 326.585 ;
      VIA 28.52 326.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 326.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 320.795 29.31 321.125 ;
      VIA 28.52 320.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 320.775 29.29 321.145 ;
      VIA 28.52 320.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 320.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 315.355 29.31 315.685 ;
      VIA 28.52 315.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 315.335 29.29 315.705 ;
      VIA 28.52 315.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 315.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 309.915 29.31 310.245 ;
      VIA 28.52 310.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 309.895 29.29 310.265 ;
      VIA 28.52 310.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 310.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 304.475 29.31 304.805 ;
      VIA 28.52 304.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 304.455 29.29 304.825 ;
      VIA 28.52 304.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 304.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 299.035 29.31 299.365 ;
      VIA 28.52 299.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 299.015 29.29 299.385 ;
      VIA 28.52 299.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 299.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 293.595 29.31 293.925 ;
      VIA 28.52 293.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 293.575 29.29 293.945 ;
      VIA 28.52 293.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 293.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 288.155 29.31 288.485 ;
      VIA 28.52 288.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 288.135 29.29 288.505 ;
      VIA 28.52 288.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 288.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 282.715 29.31 283.045 ;
      VIA 28.52 282.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 282.695 29.29 283.065 ;
      VIA 28.52 282.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 282.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 277.275 29.31 277.605 ;
      VIA 28.52 277.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 277.255 29.29 277.625 ;
      VIA 28.52 277.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 277.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 271.835 29.31 272.165 ;
      VIA 28.52 272 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 271.815 29.29 272.185 ;
      VIA 28.52 272 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 272 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 266.395 29.31 266.725 ;
      VIA 28.52 266.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 266.375 29.29 266.745 ;
      VIA 28.52 266.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 266.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 260.955 29.31 261.285 ;
      VIA 28.52 261.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 260.935 29.29 261.305 ;
      VIA 28.52 261.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 261.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 255.515 29.31 255.845 ;
      VIA 28.52 255.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 255.495 29.29 255.865 ;
      VIA 28.52 255.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 255.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 250.075 29.31 250.405 ;
      VIA 28.52 250.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 250.055 29.29 250.425 ;
      VIA 28.52 250.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 250.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 244.635 29.31 244.965 ;
      VIA 28.52 244.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 244.615 29.29 244.985 ;
      VIA 28.52 244.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 244.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 239.195 29.31 239.525 ;
      VIA 28.52 239.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 239.175 29.29 239.545 ;
      VIA 28.52 239.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 239.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 233.755 29.31 234.085 ;
      VIA 28.52 233.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 233.735 29.29 234.105 ;
      VIA 28.52 233.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 233.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 228.315 29.31 228.645 ;
      VIA 28.52 228.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 228.295 29.29 228.665 ;
      VIA 28.52 228.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 228.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 222.875 29.31 223.205 ;
      VIA 28.52 223.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 222.855 29.29 223.225 ;
      VIA 28.52 223.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 223.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 217.435 29.31 217.765 ;
      VIA 28.52 217.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 217.415 29.29 217.785 ;
      VIA 28.52 217.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 217.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 211.995 29.31 212.325 ;
      VIA 28.52 212.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 211.975 29.29 212.345 ;
      VIA 28.52 212.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 212.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 206.555 29.31 206.885 ;
      VIA 28.52 206.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 206.535 29.29 206.905 ;
      VIA 28.52 206.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 206.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 201.115 29.31 201.445 ;
      VIA 28.52 201.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 201.095 29.29 201.465 ;
      VIA 28.52 201.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 201.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 195.675 29.31 196.005 ;
      VIA 28.52 195.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 195.655 29.29 196.025 ;
      VIA 28.52 195.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 195.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 190.235 29.31 190.565 ;
      VIA 28.52 190.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 190.215 29.29 190.585 ;
      VIA 28.52 190.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 190.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 184.795 29.31 185.125 ;
      VIA 28.52 184.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 184.775 29.29 185.145 ;
      VIA 28.52 184.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 184.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 179.355 29.31 179.685 ;
      VIA 28.52 179.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 179.335 29.29 179.705 ;
      VIA 28.52 179.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 179.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 173.915 29.31 174.245 ;
      VIA 28.52 174.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 173.895 29.29 174.265 ;
      VIA 28.52 174.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 174.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 168.475 29.31 168.805 ;
      VIA 28.52 168.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 168.455 29.29 168.825 ;
      VIA 28.52 168.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 168.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 163.035 29.31 163.365 ;
      VIA 28.52 163.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 163.015 29.29 163.385 ;
      VIA 28.52 163.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 163.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 157.595 29.31 157.925 ;
      VIA 28.52 157.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 157.575 29.29 157.945 ;
      VIA 28.52 157.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 157.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 152.155 29.31 152.485 ;
      VIA 28.52 152.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 152.135 29.29 152.505 ;
      VIA 28.52 152.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 152.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 146.715 29.31 147.045 ;
      VIA 28.52 146.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 146.695 29.29 147.065 ;
      VIA 28.52 146.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 146.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 141.275 29.31 141.605 ;
      VIA 28.52 141.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 141.255 29.29 141.625 ;
      VIA 28.52 141.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 141.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 135.835 29.31 136.165 ;
      VIA 28.52 136 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 135.815 29.29 136.185 ;
      VIA 28.52 136 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 136 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 130.395 29.31 130.725 ;
      VIA 28.52 130.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 130.375 29.29 130.745 ;
      VIA 28.52 130.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 130.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 124.955 29.31 125.285 ;
      VIA 28.52 125.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 124.935 29.29 125.305 ;
      VIA 28.52 125.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 125.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 119.515 29.31 119.845 ;
      VIA 28.52 119.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 119.495 29.29 119.865 ;
      VIA 28.52 119.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 119.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 114.075 29.31 114.405 ;
      VIA 28.52 114.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 114.055 29.29 114.425 ;
      VIA 28.52 114.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 114.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 108.635 29.31 108.965 ;
      VIA 28.52 108.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 108.615 29.29 108.985 ;
      VIA 28.52 108.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 108.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 103.195 29.31 103.525 ;
      VIA 28.52 103.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 103.175 29.29 103.545 ;
      VIA 28.52 103.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 103.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 97.755 29.31 98.085 ;
      VIA 28.52 97.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 97.735 29.29 98.105 ;
      VIA 28.52 97.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 97.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 92.315 29.31 92.645 ;
      VIA 28.52 92.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 92.295 29.29 92.665 ;
      VIA 28.52 92.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 92.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 86.875 29.31 87.205 ;
      VIA 28.52 87.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 86.855 29.29 87.225 ;
      VIA 28.52 87.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 87.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 81.435 29.31 81.765 ;
      VIA 28.52 81.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 81.415 29.29 81.785 ;
      VIA 28.52 81.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 81.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 75.995 29.31 76.325 ;
      VIA 28.52 76.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 75.975 29.29 76.345 ;
      VIA 28.52 76.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 76.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 70.555 29.31 70.885 ;
      VIA 28.52 70.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 70.535 29.29 70.905 ;
      VIA 28.52 70.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 70.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 65.115 29.31 65.445 ;
      VIA 28.52 65.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 65.095 29.29 65.465 ;
      VIA 28.52 65.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 65.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 59.675 29.31 60.005 ;
      VIA 28.52 59.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 59.655 29.29 60.025 ;
      VIA 28.52 59.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 59.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 54.235 29.31 54.565 ;
      VIA 28.52 54.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 54.215 29.29 54.585 ;
      VIA 28.52 54.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 54.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 48.795 29.31 49.125 ;
      VIA 28.52 48.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 48.775 29.29 49.145 ;
      VIA 28.52 48.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 48.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 43.355 29.31 43.685 ;
      VIA 28.52 43.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 43.335 29.29 43.705 ;
      VIA 28.52 43.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 43.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 37.915 29.31 38.245 ;
      VIA 28.52 38.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 37.895 29.29 38.265 ;
      VIA 28.52 38.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 38.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 32.475 29.31 32.805 ;
      VIA 28.52 32.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 32.455 29.29 32.825 ;
      VIA 28.52 32.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 32.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 27.035 29.31 27.365 ;
      VIA 28.52 27.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 27.015 29.29 27.385 ;
      VIA 28.52 27.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 27.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 21.595 29.31 21.925 ;
      VIA 28.52 21.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 21.575 29.29 21.945 ;
      VIA 28.52 21.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 21.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 16.155 29.31 16.485 ;
      VIA 28.52 16.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 16.135 29.29 16.505 ;
      VIA 28.52 16.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 16.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 10.715 29.31 11.045 ;
      VIA 28.52 10.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 10.695 29.29 11.065 ;
      VIA 28.52 10.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 10.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  27.73 5.275 29.31 5.605 ;
      VIA 28.52 5.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  27.75 5.255 29.29 5.625 ;
      VIA 28.52 5.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 28.52 5.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      LAYER met5 ;
        RECT  14.15 695.52 151.45 697.12 ;
        RECT  14.15 668.32 151.45 669.92 ;
        RECT  14.15 641.12 151.45 642.72 ;
        RECT  14.15 613.92 151.45 615.52 ;
        RECT  14.15 586.72 151.45 588.32 ;
        RECT  14.15 559.52 151.45 561.12 ;
        RECT  14.15 532.32 151.45 533.92 ;
        RECT  14.15 505.12 151.45 506.72 ;
        RECT  14.15 477.92 151.45 479.52 ;
        RECT  14.15 450.72 151.45 452.32 ;
        RECT  14.15 423.52 151.45 425.12 ;
        RECT  14.15 396.32 151.45 397.92 ;
        RECT  14.15 369.12 151.45 370.72 ;
        RECT  14.15 341.92 151.45 343.52 ;
        RECT  14.15 314.72 151.45 316.32 ;
        RECT  14.15 287.52 151.45 289.12 ;
        RECT  14.15 260.32 151.45 261.92 ;
        RECT  14.15 233.12 151.45 234.72 ;
        RECT  14.15 205.92 151.45 207.52 ;
        RECT  14.15 178.72 151.45 180.32 ;
        RECT  14.15 151.52 151.45 153.12 ;
        RECT  14.15 124.32 151.45 125.92 ;
        RECT  14.15 97.12 151.45 98.72 ;
        RECT  14.15 69.92 151.45 71.52 ;
        RECT  14.15 42.72 151.45 44.32 ;
        RECT  14.15 15.52 151.45 17.12 ;
      LAYER met4 ;
        RECT  149.85 2.48 151.45 699.28 ;
        RECT  122.71 2.48 124.31 699.28 ;
        RECT  95.57 2.48 97.17 699.28 ;
        RECT  68.43 2.48 70.03 699.28 ;
        RECT  41.29 2.48 42.89 699.28 ;
        RECT  14.15 2.48 15.75 699.28 ;
      LAYER met1 ;
        RECT  1.38 698.8 176.18 699.28 ;
        RECT  1.38 693.36 176.18 693.84 ;
        RECT  1.38 687.92 176.18 688.4 ;
        RECT  1.38 682.48 176.18 682.96 ;
        RECT  1.38 677.04 176.18 677.52 ;
        RECT  1.38 671.6 176.18 672.08 ;
        RECT  1.38 666.16 176.18 666.64 ;
        RECT  1.38 660.72 176.18 661.2 ;
        RECT  1.38 655.28 176.18 655.76 ;
        RECT  1.38 649.84 176.18 650.32 ;
        RECT  1.38 644.4 176.18 644.88 ;
        RECT  1.38 638.96 176.18 639.44 ;
        RECT  1.38 633.52 176.18 634 ;
        RECT  1.38 628.08 176.18 628.56 ;
        RECT  1.38 622.64 176.18 623.12 ;
        RECT  1.38 617.2 176.18 617.68 ;
        RECT  1.38 611.76 176.18 612.24 ;
        RECT  1.38 606.32 176.18 606.8 ;
        RECT  1.38 600.88 176.18 601.36 ;
        RECT  1.38 595.44 176.18 595.92 ;
        RECT  1.38 590 176.18 590.48 ;
        RECT  1.38 584.56 176.18 585.04 ;
        RECT  1.38 579.12 176.18 579.6 ;
        RECT  1.38 573.68 176.18 574.16 ;
        RECT  1.38 568.24 176.18 568.72 ;
        RECT  1.38 562.8 176.18 563.28 ;
        RECT  1.38 557.36 176.18 557.84 ;
        RECT  1.38 551.92 176.18 552.4 ;
        RECT  1.38 546.48 176.18 546.96 ;
        RECT  1.38 541.04 176.18 541.52 ;
        RECT  1.38 535.6 176.18 536.08 ;
        RECT  1.38 530.16 176.18 530.64 ;
        RECT  1.38 524.72 176.18 525.2 ;
        RECT  1.38 519.28 176.18 519.76 ;
        RECT  1.38 513.84 176.18 514.32 ;
        RECT  1.38 508.4 176.18 508.88 ;
        RECT  1.38 502.96 176.18 503.44 ;
        RECT  1.38 497.52 176.18 498 ;
        RECT  1.38 492.08 176.18 492.56 ;
        RECT  1.38 486.64 176.18 487.12 ;
        RECT  1.38 481.2 176.18 481.68 ;
        RECT  1.38 475.76 176.18 476.24 ;
        RECT  1.38 470.32 176.18 470.8 ;
        RECT  1.38 464.88 176.18 465.36 ;
        RECT  1.38 459.44 176.18 459.92 ;
        RECT  1.38 454 176.18 454.48 ;
        RECT  1.38 448.56 176.18 449.04 ;
        RECT  1.38 443.12 176.18 443.6 ;
        RECT  1.38 437.68 176.18 438.16 ;
        RECT  1.38 432.24 176.18 432.72 ;
        RECT  1.38 426.8 176.18 427.28 ;
        RECT  1.38 421.36 176.18 421.84 ;
        RECT  1.38 415.92 176.18 416.4 ;
        RECT  1.38 410.48 176.18 410.96 ;
        RECT  1.38 405.04 176.18 405.52 ;
        RECT  1.38 399.6 176.18 400.08 ;
        RECT  1.38 394.16 176.18 394.64 ;
        RECT  1.38 388.72 176.18 389.2 ;
        RECT  1.38 383.28 176.18 383.76 ;
        RECT  1.38 377.84 176.18 378.32 ;
        RECT  1.38 372.4 176.18 372.88 ;
        RECT  1.38 366.96 176.18 367.44 ;
        RECT  1.38 361.52 176.18 362 ;
        RECT  1.38 356.08 176.18 356.56 ;
        RECT  1.38 350.64 176.18 351.12 ;
        RECT  1.38 345.2 176.18 345.68 ;
        RECT  1.38 339.76 176.18 340.24 ;
        RECT  1.38 334.32 176.18 334.8 ;
        RECT  1.38 328.88 176.18 329.36 ;
        RECT  1.38 323.44 176.18 323.92 ;
        RECT  1.38 318 176.18 318.48 ;
        RECT  1.38 312.56 176.18 313.04 ;
        RECT  1.38 307.12 176.18 307.6 ;
        RECT  1.38 301.68 176.18 302.16 ;
        RECT  1.38 296.24 176.18 296.72 ;
        RECT  1.38 290.8 176.18 291.28 ;
        RECT  1.38 285.36 176.18 285.84 ;
        RECT  1.38 279.92 176.18 280.4 ;
        RECT  1.38 274.48 176.18 274.96 ;
        RECT  1.38 269.04 176.18 269.52 ;
        RECT  1.38 263.6 176.18 264.08 ;
        RECT  1.38 258.16 176.18 258.64 ;
        RECT  1.38 252.72 176.18 253.2 ;
        RECT  1.38 247.28 176.18 247.76 ;
        RECT  1.38 241.84 176.18 242.32 ;
        RECT  1.38 236.4 176.18 236.88 ;
        RECT  1.38 230.96 176.18 231.44 ;
        RECT  1.38 225.52 176.18 226 ;
        RECT  1.38 220.08 176.18 220.56 ;
        RECT  1.38 214.64 176.18 215.12 ;
        RECT  1.38 209.2 176.18 209.68 ;
        RECT  1.38 203.76 176.18 204.24 ;
        RECT  1.38 198.32 176.18 198.8 ;
        RECT  1.38 192.88 176.18 193.36 ;
        RECT  1.38 187.44 176.18 187.92 ;
        RECT  1.38 182 176.18 182.48 ;
        RECT  1.38 176.56 176.18 177.04 ;
        RECT  1.38 171.12 176.18 171.6 ;
        RECT  1.38 165.68 176.18 166.16 ;
        RECT  1.38 160.24 176.18 160.72 ;
        RECT  1.38 154.8 176.18 155.28 ;
        RECT  1.38 149.36 176.18 149.84 ;
        RECT  1.38 143.92 176.18 144.4 ;
        RECT  1.38 138.48 176.18 138.96 ;
        RECT  1.38 133.04 176.18 133.52 ;
        RECT  1.38 127.6 176.18 128.08 ;
        RECT  1.38 122.16 176.18 122.64 ;
        RECT  1.38 116.72 176.18 117.2 ;
        RECT  1.38 111.28 176.18 111.76 ;
        RECT  1.38 105.84 176.18 106.32 ;
        RECT  1.38 100.4 176.18 100.88 ;
        RECT  1.38 94.96 176.18 95.44 ;
        RECT  1.38 89.52 176.18 90 ;
        RECT  1.38 84.08 176.18 84.56 ;
        RECT  1.38 78.64 176.18 79.12 ;
        RECT  1.38 73.2 176.18 73.68 ;
        RECT  1.38 67.76 176.18 68.24 ;
        RECT  1.38 62.32 176.18 62.8 ;
        RECT  1.38 56.88 176.18 57.36 ;
        RECT  1.38 51.44 176.18 51.92 ;
        RECT  1.38 46 176.18 46.48 ;
        RECT  1.38 40.56 176.18 41.04 ;
        RECT  1.38 35.12 176.18 35.6 ;
        RECT  1.38 29.68 176.18 30.16 ;
        RECT  1.38 24.24 176.18 24.72 ;
        RECT  1.38 18.8 176.18 19.28 ;
        RECT  1.38 13.36 176.18 13.84 ;
        RECT  1.38 7.92 176.18 8.4 ;
        RECT  1.38 2.48 176.18 2.96 ;
      VIA 150.65 696.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 669.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 641.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 614.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 587.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 560.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 533.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 505.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 478.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 451.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 424.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 397.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 369.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 342.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 315.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 288.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 261.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 233.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 206.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 179.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 152.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 125.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 97.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 70.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 43.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 150.65 16.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 696.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 669.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 641.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 614.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 587.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 560.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 533.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 505.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 478.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 451.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 424.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 397.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 369.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 342.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 315.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 288.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 261.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 233.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 206.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 179.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 152.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 125.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 97.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 70.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 43.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 123.51 16.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 696.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 669.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 641.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 614.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 587.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 560.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 533.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 505.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 478.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 451.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 424.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 397.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 369.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 342.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 315.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 288.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 261.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 233.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 206.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 179.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 152.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 125.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 97.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 70.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 43.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 96.37 16.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 696.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 669.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 641.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 614.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 587.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 560.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 533.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 505.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 478.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 451.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 424.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 397.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 369.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 342.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 315.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 288.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 261.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 233.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 206.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 179.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 152.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 125.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 97.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 70.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 43.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 69.23 16.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 696.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 669.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 641.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 614.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 587.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 560.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 533.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 505.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 478.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 451.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 424.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 397.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 369.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 342.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 315.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 288.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 261.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 233.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 206.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 179.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 152.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 125.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 97.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 70.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 43.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 42.09 16.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 696.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 669.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 641.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 614.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 587.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 560.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 533.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 505.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 478.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 451.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 424.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 397.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 369.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 342.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 315.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 288.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 261.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 233.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 206.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 179.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 152.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 125.12 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 97.92 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 70.72 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 43.52 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      VIA 14.95 16.32 ibex_id_stage_via5_6_1600_1600_1_1_1600_1600 ;
      LAYER met3 ;
        RECT  149.86 698.875 151.44 699.205 ;
      VIA 150.65 699.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 698.855 151.42 699.225 ;
      VIA 150.65 699.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 699.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 693.435 151.44 693.765 ;
      VIA 150.65 693.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 693.415 151.42 693.785 ;
      VIA 150.65 693.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 693.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 687.995 151.44 688.325 ;
      VIA 150.65 688.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 687.975 151.42 688.345 ;
      VIA 150.65 688.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 688.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 682.555 151.44 682.885 ;
      VIA 150.65 682.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 682.535 151.42 682.905 ;
      VIA 150.65 682.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 682.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 677.115 151.44 677.445 ;
      VIA 150.65 677.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 677.095 151.42 677.465 ;
      VIA 150.65 677.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 677.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 671.675 151.44 672.005 ;
      VIA 150.65 671.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 671.655 151.42 672.025 ;
      VIA 150.65 671.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 671.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 666.235 151.44 666.565 ;
      VIA 150.65 666.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 666.215 151.42 666.585 ;
      VIA 150.65 666.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 666.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 660.795 151.44 661.125 ;
      VIA 150.65 660.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 660.775 151.42 661.145 ;
      VIA 150.65 660.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 660.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 655.355 151.44 655.685 ;
      VIA 150.65 655.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 655.335 151.42 655.705 ;
      VIA 150.65 655.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 655.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 649.915 151.44 650.245 ;
      VIA 150.65 650.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 649.895 151.42 650.265 ;
      VIA 150.65 650.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 650.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 644.475 151.44 644.805 ;
      VIA 150.65 644.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 644.455 151.42 644.825 ;
      VIA 150.65 644.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 644.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 639.035 151.44 639.365 ;
      VIA 150.65 639.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 639.015 151.42 639.385 ;
      VIA 150.65 639.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 639.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 633.595 151.44 633.925 ;
      VIA 150.65 633.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 633.575 151.42 633.945 ;
      VIA 150.65 633.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 633.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 628.155 151.44 628.485 ;
      VIA 150.65 628.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 628.135 151.42 628.505 ;
      VIA 150.65 628.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 628.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 622.715 151.44 623.045 ;
      VIA 150.65 622.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 622.695 151.42 623.065 ;
      VIA 150.65 622.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 622.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 617.275 151.44 617.605 ;
      VIA 150.65 617.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 617.255 151.42 617.625 ;
      VIA 150.65 617.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 617.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 611.835 151.44 612.165 ;
      VIA 150.65 612 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 611.815 151.42 612.185 ;
      VIA 150.65 612 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 612 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 606.395 151.44 606.725 ;
      VIA 150.65 606.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 606.375 151.42 606.745 ;
      VIA 150.65 606.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 606.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 600.955 151.44 601.285 ;
      VIA 150.65 601.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 600.935 151.42 601.305 ;
      VIA 150.65 601.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 601.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 595.515 151.44 595.845 ;
      VIA 150.65 595.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 595.495 151.42 595.865 ;
      VIA 150.65 595.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 595.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 590.075 151.44 590.405 ;
      VIA 150.65 590.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 590.055 151.42 590.425 ;
      VIA 150.65 590.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 590.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 584.635 151.44 584.965 ;
      VIA 150.65 584.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 584.615 151.42 584.985 ;
      VIA 150.65 584.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 584.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 579.195 151.44 579.525 ;
      VIA 150.65 579.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 579.175 151.42 579.545 ;
      VIA 150.65 579.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 579.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 573.755 151.44 574.085 ;
      VIA 150.65 573.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 573.735 151.42 574.105 ;
      VIA 150.65 573.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 573.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 568.315 151.44 568.645 ;
      VIA 150.65 568.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 568.295 151.42 568.665 ;
      VIA 150.65 568.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 568.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 562.875 151.44 563.205 ;
      VIA 150.65 563.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 562.855 151.42 563.225 ;
      VIA 150.65 563.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 563.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 557.435 151.44 557.765 ;
      VIA 150.65 557.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 557.415 151.42 557.785 ;
      VIA 150.65 557.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 557.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 551.995 151.44 552.325 ;
      VIA 150.65 552.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 551.975 151.42 552.345 ;
      VIA 150.65 552.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 552.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 546.555 151.44 546.885 ;
      VIA 150.65 546.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 546.535 151.42 546.905 ;
      VIA 150.65 546.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 546.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 541.115 151.44 541.445 ;
      VIA 150.65 541.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 541.095 151.42 541.465 ;
      VIA 150.65 541.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 541.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 535.675 151.44 536.005 ;
      VIA 150.65 535.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 535.655 151.42 536.025 ;
      VIA 150.65 535.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 535.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 530.235 151.44 530.565 ;
      VIA 150.65 530.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 530.215 151.42 530.585 ;
      VIA 150.65 530.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 530.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 524.795 151.44 525.125 ;
      VIA 150.65 524.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 524.775 151.42 525.145 ;
      VIA 150.65 524.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 524.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 519.355 151.44 519.685 ;
      VIA 150.65 519.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 519.335 151.42 519.705 ;
      VIA 150.65 519.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 519.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 513.915 151.44 514.245 ;
      VIA 150.65 514.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 513.895 151.42 514.265 ;
      VIA 150.65 514.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 514.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 508.475 151.44 508.805 ;
      VIA 150.65 508.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 508.455 151.42 508.825 ;
      VIA 150.65 508.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 508.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 503.035 151.44 503.365 ;
      VIA 150.65 503.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 503.015 151.42 503.385 ;
      VIA 150.65 503.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 503.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 497.595 151.44 497.925 ;
      VIA 150.65 497.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 497.575 151.42 497.945 ;
      VIA 150.65 497.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 497.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 492.155 151.44 492.485 ;
      VIA 150.65 492.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 492.135 151.42 492.505 ;
      VIA 150.65 492.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 492.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 486.715 151.44 487.045 ;
      VIA 150.65 486.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 486.695 151.42 487.065 ;
      VIA 150.65 486.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 486.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 481.275 151.44 481.605 ;
      VIA 150.65 481.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 481.255 151.42 481.625 ;
      VIA 150.65 481.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 481.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 475.835 151.44 476.165 ;
      VIA 150.65 476 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 475.815 151.42 476.185 ;
      VIA 150.65 476 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 476 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 470.395 151.44 470.725 ;
      VIA 150.65 470.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 470.375 151.42 470.745 ;
      VIA 150.65 470.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 470.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 464.955 151.44 465.285 ;
      VIA 150.65 465.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 464.935 151.42 465.305 ;
      VIA 150.65 465.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 465.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 459.515 151.44 459.845 ;
      VIA 150.65 459.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 459.495 151.42 459.865 ;
      VIA 150.65 459.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 459.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 454.075 151.44 454.405 ;
      VIA 150.65 454.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 454.055 151.42 454.425 ;
      VIA 150.65 454.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 454.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 448.635 151.44 448.965 ;
      VIA 150.65 448.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 448.615 151.42 448.985 ;
      VIA 150.65 448.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 448.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 443.195 151.44 443.525 ;
      VIA 150.65 443.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 443.175 151.42 443.545 ;
      VIA 150.65 443.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 443.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 437.755 151.44 438.085 ;
      VIA 150.65 437.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 437.735 151.42 438.105 ;
      VIA 150.65 437.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 437.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 432.315 151.44 432.645 ;
      VIA 150.65 432.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 432.295 151.42 432.665 ;
      VIA 150.65 432.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 432.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 426.875 151.44 427.205 ;
      VIA 150.65 427.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 426.855 151.42 427.225 ;
      VIA 150.65 427.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 427.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 421.435 151.44 421.765 ;
      VIA 150.65 421.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 421.415 151.42 421.785 ;
      VIA 150.65 421.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 421.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 415.995 151.44 416.325 ;
      VIA 150.65 416.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 415.975 151.42 416.345 ;
      VIA 150.65 416.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 416.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 410.555 151.44 410.885 ;
      VIA 150.65 410.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 410.535 151.42 410.905 ;
      VIA 150.65 410.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 410.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 405.115 151.44 405.445 ;
      VIA 150.65 405.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 405.095 151.42 405.465 ;
      VIA 150.65 405.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 405.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 399.675 151.44 400.005 ;
      VIA 150.65 399.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 399.655 151.42 400.025 ;
      VIA 150.65 399.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 399.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 394.235 151.44 394.565 ;
      VIA 150.65 394.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 394.215 151.42 394.585 ;
      VIA 150.65 394.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 394.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 388.795 151.44 389.125 ;
      VIA 150.65 388.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 388.775 151.42 389.145 ;
      VIA 150.65 388.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 388.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 383.355 151.44 383.685 ;
      VIA 150.65 383.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 383.335 151.42 383.705 ;
      VIA 150.65 383.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 383.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 377.915 151.44 378.245 ;
      VIA 150.65 378.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 377.895 151.42 378.265 ;
      VIA 150.65 378.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 378.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 372.475 151.44 372.805 ;
      VIA 150.65 372.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 372.455 151.42 372.825 ;
      VIA 150.65 372.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 372.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 367.035 151.44 367.365 ;
      VIA 150.65 367.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 367.015 151.42 367.385 ;
      VIA 150.65 367.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 367.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 361.595 151.44 361.925 ;
      VIA 150.65 361.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 361.575 151.42 361.945 ;
      VIA 150.65 361.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 361.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 356.155 151.44 356.485 ;
      VIA 150.65 356.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 356.135 151.42 356.505 ;
      VIA 150.65 356.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 356.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 350.715 151.44 351.045 ;
      VIA 150.65 350.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 350.695 151.42 351.065 ;
      VIA 150.65 350.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 350.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 345.275 151.44 345.605 ;
      VIA 150.65 345.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 345.255 151.42 345.625 ;
      VIA 150.65 345.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 345.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 339.835 151.44 340.165 ;
      VIA 150.65 340 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 339.815 151.42 340.185 ;
      VIA 150.65 340 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 340 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 334.395 151.44 334.725 ;
      VIA 150.65 334.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 334.375 151.42 334.745 ;
      VIA 150.65 334.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 334.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 328.955 151.44 329.285 ;
      VIA 150.65 329.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 328.935 151.42 329.305 ;
      VIA 150.65 329.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 329.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 323.515 151.44 323.845 ;
      VIA 150.65 323.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 323.495 151.42 323.865 ;
      VIA 150.65 323.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 323.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 318.075 151.44 318.405 ;
      VIA 150.65 318.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 318.055 151.42 318.425 ;
      VIA 150.65 318.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 318.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 312.635 151.44 312.965 ;
      VIA 150.65 312.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 312.615 151.42 312.985 ;
      VIA 150.65 312.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 312.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 307.195 151.44 307.525 ;
      VIA 150.65 307.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 307.175 151.42 307.545 ;
      VIA 150.65 307.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 307.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 301.755 151.44 302.085 ;
      VIA 150.65 301.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 301.735 151.42 302.105 ;
      VIA 150.65 301.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 301.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 296.315 151.44 296.645 ;
      VIA 150.65 296.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 296.295 151.42 296.665 ;
      VIA 150.65 296.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 296.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 290.875 151.44 291.205 ;
      VIA 150.65 291.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 290.855 151.42 291.225 ;
      VIA 150.65 291.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 291.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 285.435 151.44 285.765 ;
      VIA 150.65 285.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 285.415 151.42 285.785 ;
      VIA 150.65 285.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 285.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 279.995 151.44 280.325 ;
      VIA 150.65 280.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 279.975 151.42 280.345 ;
      VIA 150.65 280.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 280.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 274.555 151.44 274.885 ;
      VIA 150.65 274.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 274.535 151.42 274.905 ;
      VIA 150.65 274.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 274.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 269.115 151.44 269.445 ;
      VIA 150.65 269.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 269.095 151.42 269.465 ;
      VIA 150.65 269.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 269.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 263.675 151.44 264.005 ;
      VIA 150.65 263.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 263.655 151.42 264.025 ;
      VIA 150.65 263.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 263.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 258.235 151.44 258.565 ;
      VIA 150.65 258.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 258.215 151.42 258.585 ;
      VIA 150.65 258.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 258.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 252.795 151.44 253.125 ;
      VIA 150.65 252.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 252.775 151.42 253.145 ;
      VIA 150.65 252.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 252.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 247.355 151.44 247.685 ;
      VIA 150.65 247.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 247.335 151.42 247.705 ;
      VIA 150.65 247.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 247.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 241.915 151.44 242.245 ;
      VIA 150.65 242.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 241.895 151.42 242.265 ;
      VIA 150.65 242.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 242.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 236.475 151.44 236.805 ;
      VIA 150.65 236.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 236.455 151.42 236.825 ;
      VIA 150.65 236.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 236.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 231.035 151.44 231.365 ;
      VIA 150.65 231.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 231.015 151.42 231.385 ;
      VIA 150.65 231.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 231.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 225.595 151.44 225.925 ;
      VIA 150.65 225.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 225.575 151.42 225.945 ;
      VIA 150.65 225.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 225.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 220.155 151.44 220.485 ;
      VIA 150.65 220.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 220.135 151.42 220.505 ;
      VIA 150.65 220.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 220.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 214.715 151.44 215.045 ;
      VIA 150.65 214.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 214.695 151.42 215.065 ;
      VIA 150.65 214.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 214.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 209.275 151.44 209.605 ;
      VIA 150.65 209.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 209.255 151.42 209.625 ;
      VIA 150.65 209.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 209.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 203.835 151.44 204.165 ;
      VIA 150.65 204 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 203.815 151.42 204.185 ;
      VIA 150.65 204 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 204 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 198.395 151.44 198.725 ;
      VIA 150.65 198.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 198.375 151.42 198.745 ;
      VIA 150.65 198.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 198.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 192.955 151.44 193.285 ;
      VIA 150.65 193.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 192.935 151.42 193.305 ;
      VIA 150.65 193.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 193.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 187.515 151.44 187.845 ;
      VIA 150.65 187.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 187.495 151.42 187.865 ;
      VIA 150.65 187.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 187.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 182.075 151.44 182.405 ;
      VIA 150.65 182.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 182.055 151.42 182.425 ;
      VIA 150.65 182.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 182.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 176.635 151.44 176.965 ;
      VIA 150.65 176.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 176.615 151.42 176.985 ;
      VIA 150.65 176.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 176.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 171.195 151.44 171.525 ;
      VIA 150.65 171.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 171.175 151.42 171.545 ;
      VIA 150.65 171.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 171.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 165.755 151.44 166.085 ;
      VIA 150.65 165.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 165.735 151.42 166.105 ;
      VIA 150.65 165.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 165.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 160.315 151.44 160.645 ;
      VIA 150.65 160.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 160.295 151.42 160.665 ;
      VIA 150.65 160.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 160.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 154.875 151.44 155.205 ;
      VIA 150.65 155.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 154.855 151.42 155.225 ;
      VIA 150.65 155.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 155.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 149.435 151.44 149.765 ;
      VIA 150.65 149.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 149.415 151.42 149.785 ;
      VIA 150.65 149.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 149.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 143.995 151.44 144.325 ;
      VIA 150.65 144.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 143.975 151.42 144.345 ;
      VIA 150.65 144.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 144.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 138.555 151.44 138.885 ;
      VIA 150.65 138.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 138.535 151.42 138.905 ;
      VIA 150.65 138.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 138.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 133.115 151.44 133.445 ;
      VIA 150.65 133.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 133.095 151.42 133.465 ;
      VIA 150.65 133.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 133.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 127.675 151.44 128.005 ;
      VIA 150.65 127.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 127.655 151.42 128.025 ;
      VIA 150.65 127.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 127.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 122.235 151.44 122.565 ;
      VIA 150.65 122.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 122.215 151.42 122.585 ;
      VIA 150.65 122.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 122.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 116.795 151.44 117.125 ;
      VIA 150.65 116.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 116.775 151.42 117.145 ;
      VIA 150.65 116.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 116.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 111.355 151.44 111.685 ;
      VIA 150.65 111.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 111.335 151.42 111.705 ;
      VIA 150.65 111.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 111.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 105.915 151.44 106.245 ;
      VIA 150.65 106.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 105.895 151.42 106.265 ;
      VIA 150.65 106.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 106.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 100.475 151.44 100.805 ;
      VIA 150.65 100.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 100.455 151.42 100.825 ;
      VIA 150.65 100.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 100.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 95.035 151.44 95.365 ;
      VIA 150.65 95.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 95.015 151.42 95.385 ;
      VIA 150.65 95.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 95.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 89.595 151.44 89.925 ;
      VIA 150.65 89.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 89.575 151.42 89.945 ;
      VIA 150.65 89.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 89.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 84.155 151.44 84.485 ;
      VIA 150.65 84.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 84.135 151.42 84.505 ;
      VIA 150.65 84.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 84.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 78.715 151.44 79.045 ;
      VIA 150.65 78.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 78.695 151.42 79.065 ;
      VIA 150.65 78.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 78.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 73.275 151.44 73.605 ;
      VIA 150.65 73.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 73.255 151.42 73.625 ;
      VIA 150.65 73.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 73.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 67.835 151.44 68.165 ;
      VIA 150.65 68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 67.815 151.42 68.185 ;
      VIA 150.65 68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 62.395 151.44 62.725 ;
      VIA 150.65 62.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 62.375 151.42 62.745 ;
      VIA 150.65 62.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 62.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 56.955 151.44 57.285 ;
      VIA 150.65 57.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 56.935 151.42 57.305 ;
      VIA 150.65 57.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 57.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 51.515 151.44 51.845 ;
      VIA 150.65 51.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 51.495 151.42 51.865 ;
      VIA 150.65 51.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 51.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 46.075 151.44 46.405 ;
      VIA 150.65 46.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 46.055 151.42 46.425 ;
      VIA 150.65 46.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 46.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 40.635 151.44 40.965 ;
      VIA 150.65 40.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 40.615 151.42 40.985 ;
      VIA 150.65 40.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 40.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 35.195 151.44 35.525 ;
      VIA 150.65 35.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 35.175 151.42 35.545 ;
      VIA 150.65 35.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 35.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 29.755 151.44 30.085 ;
      VIA 150.65 29.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 29.735 151.42 30.105 ;
      VIA 150.65 29.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 29.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 24.315 151.44 24.645 ;
      VIA 150.65 24.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 24.295 151.42 24.665 ;
      VIA 150.65 24.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 24.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 18.875 151.44 19.205 ;
      VIA 150.65 19.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 18.855 151.42 19.225 ;
      VIA 150.65 19.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 19.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 13.435 151.44 13.765 ;
      VIA 150.65 13.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 13.415 151.42 13.785 ;
      VIA 150.65 13.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 13.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 7.995 151.44 8.325 ;
      VIA 150.65 8.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 7.975 151.42 8.345 ;
      VIA 150.65 8.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 8.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  149.86 2.555 151.44 2.885 ;
      VIA 150.65 2.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  149.88 2.535 151.42 2.905 ;
      VIA 150.65 2.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 150.65 2.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 698.875 124.3 699.205 ;
      VIA 123.51 699.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 698.855 124.28 699.225 ;
      VIA 123.51 699.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 699.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 693.435 124.3 693.765 ;
      VIA 123.51 693.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 693.415 124.28 693.785 ;
      VIA 123.51 693.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 693.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 687.995 124.3 688.325 ;
      VIA 123.51 688.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 687.975 124.28 688.345 ;
      VIA 123.51 688.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 688.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 682.555 124.3 682.885 ;
      VIA 123.51 682.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 682.535 124.28 682.905 ;
      VIA 123.51 682.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 682.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 677.115 124.3 677.445 ;
      VIA 123.51 677.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 677.095 124.28 677.465 ;
      VIA 123.51 677.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 677.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 671.675 124.3 672.005 ;
      VIA 123.51 671.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 671.655 124.28 672.025 ;
      VIA 123.51 671.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 671.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 666.235 124.3 666.565 ;
      VIA 123.51 666.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 666.215 124.28 666.585 ;
      VIA 123.51 666.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 666.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 660.795 124.3 661.125 ;
      VIA 123.51 660.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 660.775 124.28 661.145 ;
      VIA 123.51 660.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 660.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 655.355 124.3 655.685 ;
      VIA 123.51 655.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 655.335 124.28 655.705 ;
      VIA 123.51 655.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 655.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 649.915 124.3 650.245 ;
      VIA 123.51 650.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 649.895 124.28 650.265 ;
      VIA 123.51 650.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 650.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 644.475 124.3 644.805 ;
      VIA 123.51 644.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 644.455 124.28 644.825 ;
      VIA 123.51 644.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 644.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 639.035 124.3 639.365 ;
      VIA 123.51 639.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 639.015 124.28 639.385 ;
      VIA 123.51 639.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 639.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 633.595 124.3 633.925 ;
      VIA 123.51 633.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 633.575 124.28 633.945 ;
      VIA 123.51 633.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 633.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 628.155 124.3 628.485 ;
      VIA 123.51 628.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 628.135 124.28 628.505 ;
      VIA 123.51 628.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 628.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 622.715 124.3 623.045 ;
      VIA 123.51 622.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 622.695 124.28 623.065 ;
      VIA 123.51 622.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 622.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 617.275 124.3 617.605 ;
      VIA 123.51 617.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 617.255 124.28 617.625 ;
      VIA 123.51 617.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 617.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 611.835 124.3 612.165 ;
      VIA 123.51 612 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 611.815 124.28 612.185 ;
      VIA 123.51 612 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 612 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 606.395 124.3 606.725 ;
      VIA 123.51 606.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 606.375 124.28 606.745 ;
      VIA 123.51 606.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 606.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 600.955 124.3 601.285 ;
      VIA 123.51 601.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 600.935 124.28 601.305 ;
      VIA 123.51 601.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 601.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 595.515 124.3 595.845 ;
      VIA 123.51 595.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 595.495 124.28 595.865 ;
      VIA 123.51 595.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 595.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 590.075 124.3 590.405 ;
      VIA 123.51 590.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 590.055 124.28 590.425 ;
      VIA 123.51 590.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 590.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 584.635 124.3 584.965 ;
      VIA 123.51 584.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 584.615 124.28 584.985 ;
      VIA 123.51 584.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 584.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 579.195 124.3 579.525 ;
      VIA 123.51 579.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 579.175 124.28 579.545 ;
      VIA 123.51 579.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 579.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 573.755 124.3 574.085 ;
      VIA 123.51 573.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 573.735 124.28 574.105 ;
      VIA 123.51 573.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 573.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 568.315 124.3 568.645 ;
      VIA 123.51 568.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 568.295 124.28 568.665 ;
      VIA 123.51 568.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 568.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 562.875 124.3 563.205 ;
      VIA 123.51 563.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 562.855 124.28 563.225 ;
      VIA 123.51 563.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 563.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 557.435 124.3 557.765 ;
      VIA 123.51 557.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 557.415 124.28 557.785 ;
      VIA 123.51 557.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 557.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 551.995 124.3 552.325 ;
      VIA 123.51 552.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 551.975 124.28 552.345 ;
      VIA 123.51 552.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 552.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 546.555 124.3 546.885 ;
      VIA 123.51 546.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 546.535 124.28 546.905 ;
      VIA 123.51 546.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 546.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 541.115 124.3 541.445 ;
      VIA 123.51 541.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 541.095 124.28 541.465 ;
      VIA 123.51 541.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 541.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 535.675 124.3 536.005 ;
      VIA 123.51 535.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 535.655 124.28 536.025 ;
      VIA 123.51 535.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 535.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 530.235 124.3 530.565 ;
      VIA 123.51 530.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 530.215 124.28 530.585 ;
      VIA 123.51 530.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 530.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 524.795 124.3 525.125 ;
      VIA 123.51 524.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 524.775 124.28 525.145 ;
      VIA 123.51 524.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 524.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 519.355 124.3 519.685 ;
      VIA 123.51 519.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 519.335 124.28 519.705 ;
      VIA 123.51 519.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 519.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 513.915 124.3 514.245 ;
      VIA 123.51 514.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 513.895 124.28 514.265 ;
      VIA 123.51 514.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 514.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 508.475 124.3 508.805 ;
      VIA 123.51 508.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 508.455 124.28 508.825 ;
      VIA 123.51 508.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 508.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 503.035 124.3 503.365 ;
      VIA 123.51 503.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 503.015 124.28 503.385 ;
      VIA 123.51 503.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 503.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 497.595 124.3 497.925 ;
      VIA 123.51 497.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 497.575 124.28 497.945 ;
      VIA 123.51 497.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 497.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 492.155 124.3 492.485 ;
      VIA 123.51 492.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 492.135 124.28 492.505 ;
      VIA 123.51 492.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 492.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 486.715 124.3 487.045 ;
      VIA 123.51 486.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 486.695 124.28 487.065 ;
      VIA 123.51 486.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 486.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 481.275 124.3 481.605 ;
      VIA 123.51 481.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 481.255 124.28 481.625 ;
      VIA 123.51 481.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 481.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 475.835 124.3 476.165 ;
      VIA 123.51 476 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 475.815 124.28 476.185 ;
      VIA 123.51 476 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 476 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 470.395 124.3 470.725 ;
      VIA 123.51 470.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 470.375 124.28 470.745 ;
      VIA 123.51 470.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 470.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 464.955 124.3 465.285 ;
      VIA 123.51 465.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 464.935 124.28 465.305 ;
      VIA 123.51 465.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 465.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 459.515 124.3 459.845 ;
      VIA 123.51 459.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 459.495 124.28 459.865 ;
      VIA 123.51 459.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 459.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 454.075 124.3 454.405 ;
      VIA 123.51 454.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 454.055 124.28 454.425 ;
      VIA 123.51 454.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 454.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 448.635 124.3 448.965 ;
      VIA 123.51 448.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 448.615 124.28 448.985 ;
      VIA 123.51 448.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 448.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 443.195 124.3 443.525 ;
      VIA 123.51 443.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 443.175 124.28 443.545 ;
      VIA 123.51 443.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 443.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 437.755 124.3 438.085 ;
      VIA 123.51 437.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 437.735 124.28 438.105 ;
      VIA 123.51 437.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 437.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 432.315 124.3 432.645 ;
      VIA 123.51 432.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 432.295 124.28 432.665 ;
      VIA 123.51 432.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 432.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 426.875 124.3 427.205 ;
      VIA 123.51 427.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 426.855 124.28 427.225 ;
      VIA 123.51 427.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 427.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 421.435 124.3 421.765 ;
      VIA 123.51 421.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 421.415 124.28 421.785 ;
      VIA 123.51 421.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 421.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 415.995 124.3 416.325 ;
      VIA 123.51 416.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 415.975 124.28 416.345 ;
      VIA 123.51 416.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 416.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 410.555 124.3 410.885 ;
      VIA 123.51 410.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 410.535 124.28 410.905 ;
      VIA 123.51 410.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 410.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 405.115 124.3 405.445 ;
      VIA 123.51 405.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 405.095 124.28 405.465 ;
      VIA 123.51 405.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 405.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 399.675 124.3 400.005 ;
      VIA 123.51 399.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 399.655 124.28 400.025 ;
      VIA 123.51 399.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 399.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 394.235 124.3 394.565 ;
      VIA 123.51 394.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 394.215 124.28 394.585 ;
      VIA 123.51 394.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 394.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 388.795 124.3 389.125 ;
      VIA 123.51 388.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 388.775 124.28 389.145 ;
      VIA 123.51 388.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 388.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 383.355 124.3 383.685 ;
      VIA 123.51 383.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 383.335 124.28 383.705 ;
      VIA 123.51 383.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 383.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 377.915 124.3 378.245 ;
      VIA 123.51 378.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 377.895 124.28 378.265 ;
      VIA 123.51 378.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 378.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 372.475 124.3 372.805 ;
      VIA 123.51 372.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 372.455 124.28 372.825 ;
      VIA 123.51 372.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 372.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 367.035 124.3 367.365 ;
      VIA 123.51 367.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 367.015 124.28 367.385 ;
      VIA 123.51 367.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 367.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 361.595 124.3 361.925 ;
      VIA 123.51 361.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 361.575 124.28 361.945 ;
      VIA 123.51 361.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 361.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 356.155 124.3 356.485 ;
      VIA 123.51 356.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 356.135 124.28 356.505 ;
      VIA 123.51 356.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 356.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 350.715 124.3 351.045 ;
      VIA 123.51 350.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 350.695 124.28 351.065 ;
      VIA 123.51 350.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 350.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 345.275 124.3 345.605 ;
      VIA 123.51 345.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 345.255 124.28 345.625 ;
      VIA 123.51 345.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 345.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 339.835 124.3 340.165 ;
      VIA 123.51 340 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 339.815 124.28 340.185 ;
      VIA 123.51 340 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 340 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 334.395 124.3 334.725 ;
      VIA 123.51 334.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 334.375 124.28 334.745 ;
      VIA 123.51 334.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 334.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 328.955 124.3 329.285 ;
      VIA 123.51 329.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 328.935 124.28 329.305 ;
      VIA 123.51 329.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 329.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 323.515 124.3 323.845 ;
      VIA 123.51 323.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 323.495 124.28 323.865 ;
      VIA 123.51 323.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 323.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 318.075 124.3 318.405 ;
      VIA 123.51 318.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 318.055 124.28 318.425 ;
      VIA 123.51 318.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 318.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 312.635 124.3 312.965 ;
      VIA 123.51 312.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 312.615 124.28 312.985 ;
      VIA 123.51 312.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 312.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 307.195 124.3 307.525 ;
      VIA 123.51 307.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 307.175 124.28 307.545 ;
      VIA 123.51 307.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 307.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 301.755 124.3 302.085 ;
      VIA 123.51 301.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 301.735 124.28 302.105 ;
      VIA 123.51 301.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 301.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 296.315 124.3 296.645 ;
      VIA 123.51 296.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 296.295 124.28 296.665 ;
      VIA 123.51 296.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 296.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 290.875 124.3 291.205 ;
      VIA 123.51 291.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 290.855 124.28 291.225 ;
      VIA 123.51 291.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 291.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 285.435 124.3 285.765 ;
      VIA 123.51 285.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 285.415 124.28 285.785 ;
      VIA 123.51 285.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 285.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 279.995 124.3 280.325 ;
      VIA 123.51 280.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 279.975 124.28 280.345 ;
      VIA 123.51 280.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 280.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 274.555 124.3 274.885 ;
      VIA 123.51 274.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 274.535 124.28 274.905 ;
      VIA 123.51 274.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 274.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 269.115 124.3 269.445 ;
      VIA 123.51 269.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 269.095 124.28 269.465 ;
      VIA 123.51 269.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 269.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 263.675 124.3 264.005 ;
      VIA 123.51 263.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 263.655 124.28 264.025 ;
      VIA 123.51 263.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 263.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 258.235 124.3 258.565 ;
      VIA 123.51 258.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 258.215 124.28 258.585 ;
      VIA 123.51 258.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 258.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 252.795 124.3 253.125 ;
      VIA 123.51 252.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 252.775 124.28 253.145 ;
      VIA 123.51 252.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 252.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 247.355 124.3 247.685 ;
      VIA 123.51 247.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 247.335 124.28 247.705 ;
      VIA 123.51 247.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 247.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 241.915 124.3 242.245 ;
      VIA 123.51 242.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 241.895 124.28 242.265 ;
      VIA 123.51 242.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 242.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 236.475 124.3 236.805 ;
      VIA 123.51 236.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 236.455 124.28 236.825 ;
      VIA 123.51 236.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 236.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 231.035 124.3 231.365 ;
      VIA 123.51 231.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 231.015 124.28 231.385 ;
      VIA 123.51 231.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 231.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 225.595 124.3 225.925 ;
      VIA 123.51 225.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 225.575 124.28 225.945 ;
      VIA 123.51 225.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 225.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 220.155 124.3 220.485 ;
      VIA 123.51 220.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 220.135 124.28 220.505 ;
      VIA 123.51 220.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 220.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 214.715 124.3 215.045 ;
      VIA 123.51 214.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 214.695 124.28 215.065 ;
      VIA 123.51 214.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 214.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 209.275 124.3 209.605 ;
      VIA 123.51 209.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 209.255 124.28 209.625 ;
      VIA 123.51 209.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 209.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 203.835 124.3 204.165 ;
      VIA 123.51 204 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 203.815 124.28 204.185 ;
      VIA 123.51 204 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 204 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 198.395 124.3 198.725 ;
      VIA 123.51 198.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 198.375 124.28 198.745 ;
      VIA 123.51 198.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 198.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 192.955 124.3 193.285 ;
      VIA 123.51 193.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 192.935 124.28 193.305 ;
      VIA 123.51 193.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 193.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 187.515 124.3 187.845 ;
      VIA 123.51 187.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 187.495 124.28 187.865 ;
      VIA 123.51 187.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 187.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 182.075 124.3 182.405 ;
      VIA 123.51 182.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 182.055 124.28 182.425 ;
      VIA 123.51 182.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 182.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 176.635 124.3 176.965 ;
      VIA 123.51 176.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 176.615 124.28 176.985 ;
      VIA 123.51 176.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 176.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 171.195 124.3 171.525 ;
      VIA 123.51 171.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 171.175 124.28 171.545 ;
      VIA 123.51 171.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 171.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 165.755 124.3 166.085 ;
      VIA 123.51 165.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 165.735 124.28 166.105 ;
      VIA 123.51 165.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 165.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 160.315 124.3 160.645 ;
      VIA 123.51 160.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 160.295 124.28 160.665 ;
      VIA 123.51 160.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 160.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 154.875 124.3 155.205 ;
      VIA 123.51 155.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 154.855 124.28 155.225 ;
      VIA 123.51 155.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 155.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 149.435 124.3 149.765 ;
      VIA 123.51 149.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 149.415 124.28 149.785 ;
      VIA 123.51 149.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 149.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 143.995 124.3 144.325 ;
      VIA 123.51 144.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 143.975 124.28 144.345 ;
      VIA 123.51 144.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 144.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 138.555 124.3 138.885 ;
      VIA 123.51 138.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 138.535 124.28 138.905 ;
      VIA 123.51 138.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 138.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 133.115 124.3 133.445 ;
      VIA 123.51 133.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 133.095 124.28 133.465 ;
      VIA 123.51 133.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 133.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 127.675 124.3 128.005 ;
      VIA 123.51 127.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 127.655 124.28 128.025 ;
      VIA 123.51 127.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 127.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 122.235 124.3 122.565 ;
      VIA 123.51 122.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 122.215 124.28 122.585 ;
      VIA 123.51 122.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 122.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 116.795 124.3 117.125 ;
      VIA 123.51 116.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 116.775 124.28 117.145 ;
      VIA 123.51 116.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 116.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 111.355 124.3 111.685 ;
      VIA 123.51 111.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 111.335 124.28 111.705 ;
      VIA 123.51 111.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 111.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 105.915 124.3 106.245 ;
      VIA 123.51 106.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 105.895 124.28 106.265 ;
      VIA 123.51 106.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 106.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 100.475 124.3 100.805 ;
      VIA 123.51 100.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 100.455 124.28 100.825 ;
      VIA 123.51 100.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 100.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 95.035 124.3 95.365 ;
      VIA 123.51 95.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 95.015 124.28 95.385 ;
      VIA 123.51 95.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 95.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 89.595 124.3 89.925 ;
      VIA 123.51 89.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 89.575 124.28 89.945 ;
      VIA 123.51 89.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 89.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 84.155 124.3 84.485 ;
      VIA 123.51 84.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 84.135 124.28 84.505 ;
      VIA 123.51 84.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 84.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 78.715 124.3 79.045 ;
      VIA 123.51 78.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 78.695 124.28 79.065 ;
      VIA 123.51 78.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 78.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 73.275 124.3 73.605 ;
      VIA 123.51 73.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 73.255 124.28 73.625 ;
      VIA 123.51 73.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 73.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 67.835 124.3 68.165 ;
      VIA 123.51 68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 67.815 124.28 68.185 ;
      VIA 123.51 68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 62.395 124.3 62.725 ;
      VIA 123.51 62.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 62.375 124.28 62.745 ;
      VIA 123.51 62.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 62.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 56.955 124.3 57.285 ;
      VIA 123.51 57.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 56.935 124.28 57.305 ;
      VIA 123.51 57.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 57.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 51.515 124.3 51.845 ;
      VIA 123.51 51.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 51.495 124.28 51.865 ;
      VIA 123.51 51.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 51.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 46.075 124.3 46.405 ;
      VIA 123.51 46.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 46.055 124.28 46.425 ;
      VIA 123.51 46.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 46.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 40.635 124.3 40.965 ;
      VIA 123.51 40.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 40.615 124.28 40.985 ;
      VIA 123.51 40.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 40.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 35.195 124.3 35.525 ;
      VIA 123.51 35.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 35.175 124.28 35.545 ;
      VIA 123.51 35.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 35.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 29.755 124.3 30.085 ;
      VIA 123.51 29.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 29.735 124.28 30.105 ;
      VIA 123.51 29.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 29.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 24.315 124.3 24.645 ;
      VIA 123.51 24.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 24.295 124.28 24.665 ;
      VIA 123.51 24.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 24.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 18.875 124.3 19.205 ;
      VIA 123.51 19.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 18.855 124.28 19.225 ;
      VIA 123.51 19.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 19.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 13.435 124.3 13.765 ;
      VIA 123.51 13.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 13.415 124.28 13.785 ;
      VIA 123.51 13.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 13.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 7.995 124.3 8.325 ;
      VIA 123.51 8.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 7.975 124.28 8.345 ;
      VIA 123.51 8.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 8.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  122.72 2.555 124.3 2.885 ;
      VIA 123.51 2.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  122.74 2.535 124.28 2.905 ;
      VIA 123.51 2.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 123.51 2.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 698.875 97.16 699.205 ;
      VIA 96.37 699.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 698.855 97.14 699.225 ;
      VIA 96.37 699.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 699.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 693.435 97.16 693.765 ;
      VIA 96.37 693.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 693.415 97.14 693.785 ;
      VIA 96.37 693.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 693.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 687.995 97.16 688.325 ;
      VIA 96.37 688.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 687.975 97.14 688.345 ;
      VIA 96.37 688.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 688.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 682.555 97.16 682.885 ;
      VIA 96.37 682.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 682.535 97.14 682.905 ;
      VIA 96.37 682.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 682.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 677.115 97.16 677.445 ;
      VIA 96.37 677.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 677.095 97.14 677.465 ;
      VIA 96.37 677.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 677.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 671.675 97.16 672.005 ;
      VIA 96.37 671.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 671.655 97.14 672.025 ;
      VIA 96.37 671.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 671.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 666.235 97.16 666.565 ;
      VIA 96.37 666.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 666.215 97.14 666.585 ;
      VIA 96.37 666.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 666.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 660.795 97.16 661.125 ;
      VIA 96.37 660.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 660.775 97.14 661.145 ;
      VIA 96.37 660.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 660.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 655.355 97.16 655.685 ;
      VIA 96.37 655.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 655.335 97.14 655.705 ;
      VIA 96.37 655.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 655.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 649.915 97.16 650.245 ;
      VIA 96.37 650.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 649.895 97.14 650.265 ;
      VIA 96.37 650.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 650.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 644.475 97.16 644.805 ;
      VIA 96.37 644.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 644.455 97.14 644.825 ;
      VIA 96.37 644.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 644.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 639.035 97.16 639.365 ;
      VIA 96.37 639.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 639.015 97.14 639.385 ;
      VIA 96.37 639.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 639.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 633.595 97.16 633.925 ;
      VIA 96.37 633.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 633.575 97.14 633.945 ;
      VIA 96.37 633.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 633.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 628.155 97.16 628.485 ;
      VIA 96.37 628.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 628.135 97.14 628.505 ;
      VIA 96.37 628.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 628.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 622.715 97.16 623.045 ;
      VIA 96.37 622.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 622.695 97.14 623.065 ;
      VIA 96.37 622.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 622.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 617.275 97.16 617.605 ;
      VIA 96.37 617.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 617.255 97.14 617.625 ;
      VIA 96.37 617.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 617.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 611.835 97.16 612.165 ;
      VIA 96.37 612 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 611.815 97.14 612.185 ;
      VIA 96.37 612 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 612 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 606.395 97.16 606.725 ;
      VIA 96.37 606.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 606.375 97.14 606.745 ;
      VIA 96.37 606.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 606.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 600.955 97.16 601.285 ;
      VIA 96.37 601.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 600.935 97.14 601.305 ;
      VIA 96.37 601.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 601.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 595.515 97.16 595.845 ;
      VIA 96.37 595.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 595.495 97.14 595.865 ;
      VIA 96.37 595.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 595.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 590.075 97.16 590.405 ;
      VIA 96.37 590.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 590.055 97.14 590.425 ;
      VIA 96.37 590.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 590.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 584.635 97.16 584.965 ;
      VIA 96.37 584.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 584.615 97.14 584.985 ;
      VIA 96.37 584.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 584.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 579.195 97.16 579.525 ;
      VIA 96.37 579.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 579.175 97.14 579.545 ;
      VIA 96.37 579.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 579.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 573.755 97.16 574.085 ;
      VIA 96.37 573.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 573.735 97.14 574.105 ;
      VIA 96.37 573.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 573.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 568.315 97.16 568.645 ;
      VIA 96.37 568.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 568.295 97.14 568.665 ;
      VIA 96.37 568.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 568.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 562.875 97.16 563.205 ;
      VIA 96.37 563.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 562.855 97.14 563.225 ;
      VIA 96.37 563.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 563.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 557.435 97.16 557.765 ;
      VIA 96.37 557.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 557.415 97.14 557.785 ;
      VIA 96.37 557.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 557.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 551.995 97.16 552.325 ;
      VIA 96.37 552.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 551.975 97.14 552.345 ;
      VIA 96.37 552.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 552.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 546.555 97.16 546.885 ;
      VIA 96.37 546.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 546.535 97.14 546.905 ;
      VIA 96.37 546.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 546.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 541.115 97.16 541.445 ;
      VIA 96.37 541.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 541.095 97.14 541.465 ;
      VIA 96.37 541.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 541.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 535.675 97.16 536.005 ;
      VIA 96.37 535.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 535.655 97.14 536.025 ;
      VIA 96.37 535.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 535.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 530.235 97.16 530.565 ;
      VIA 96.37 530.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 530.215 97.14 530.585 ;
      VIA 96.37 530.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 530.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 524.795 97.16 525.125 ;
      VIA 96.37 524.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 524.775 97.14 525.145 ;
      VIA 96.37 524.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 524.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 519.355 97.16 519.685 ;
      VIA 96.37 519.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 519.335 97.14 519.705 ;
      VIA 96.37 519.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 519.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 513.915 97.16 514.245 ;
      VIA 96.37 514.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 513.895 97.14 514.265 ;
      VIA 96.37 514.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 514.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 508.475 97.16 508.805 ;
      VIA 96.37 508.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 508.455 97.14 508.825 ;
      VIA 96.37 508.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 508.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 503.035 97.16 503.365 ;
      VIA 96.37 503.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 503.015 97.14 503.385 ;
      VIA 96.37 503.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 503.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 497.595 97.16 497.925 ;
      VIA 96.37 497.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 497.575 97.14 497.945 ;
      VIA 96.37 497.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 497.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 492.155 97.16 492.485 ;
      VIA 96.37 492.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 492.135 97.14 492.505 ;
      VIA 96.37 492.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 492.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 486.715 97.16 487.045 ;
      VIA 96.37 486.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 486.695 97.14 487.065 ;
      VIA 96.37 486.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 486.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 481.275 97.16 481.605 ;
      VIA 96.37 481.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 481.255 97.14 481.625 ;
      VIA 96.37 481.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 481.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 475.835 97.16 476.165 ;
      VIA 96.37 476 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 475.815 97.14 476.185 ;
      VIA 96.37 476 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 476 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 470.395 97.16 470.725 ;
      VIA 96.37 470.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 470.375 97.14 470.745 ;
      VIA 96.37 470.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 470.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 464.955 97.16 465.285 ;
      VIA 96.37 465.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 464.935 97.14 465.305 ;
      VIA 96.37 465.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 465.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 459.515 97.16 459.845 ;
      VIA 96.37 459.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 459.495 97.14 459.865 ;
      VIA 96.37 459.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 459.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 454.075 97.16 454.405 ;
      VIA 96.37 454.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 454.055 97.14 454.425 ;
      VIA 96.37 454.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 454.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 448.635 97.16 448.965 ;
      VIA 96.37 448.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 448.615 97.14 448.985 ;
      VIA 96.37 448.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 448.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 443.195 97.16 443.525 ;
      VIA 96.37 443.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 443.175 97.14 443.545 ;
      VIA 96.37 443.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 443.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 437.755 97.16 438.085 ;
      VIA 96.37 437.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 437.735 97.14 438.105 ;
      VIA 96.37 437.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 437.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 432.315 97.16 432.645 ;
      VIA 96.37 432.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 432.295 97.14 432.665 ;
      VIA 96.37 432.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 432.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 426.875 97.16 427.205 ;
      VIA 96.37 427.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 426.855 97.14 427.225 ;
      VIA 96.37 427.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 427.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 421.435 97.16 421.765 ;
      VIA 96.37 421.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 421.415 97.14 421.785 ;
      VIA 96.37 421.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 421.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 415.995 97.16 416.325 ;
      VIA 96.37 416.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 415.975 97.14 416.345 ;
      VIA 96.37 416.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 416.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 410.555 97.16 410.885 ;
      VIA 96.37 410.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 410.535 97.14 410.905 ;
      VIA 96.37 410.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 410.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 405.115 97.16 405.445 ;
      VIA 96.37 405.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 405.095 97.14 405.465 ;
      VIA 96.37 405.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 405.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 399.675 97.16 400.005 ;
      VIA 96.37 399.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 399.655 97.14 400.025 ;
      VIA 96.37 399.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 399.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 394.235 97.16 394.565 ;
      VIA 96.37 394.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 394.215 97.14 394.585 ;
      VIA 96.37 394.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 394.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 388.795 97.16 389.125 ;
      VIA 96.37 388.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 388.775 97.14 389.145 ;
      VIA 96.37 388.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 388.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 383.355 97.16 383.685 ;
      VIA 96.37 383.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 383.335 97.14 383.705 ;
      VIA 96.37 383.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 383.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 377.915 97.16 378.245 ;
      VIA 96.37 378.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 377.895 97.14 378.265 ;
      VIA 96.37 378.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 378.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 372.475 97.16 372.805 ;
      VIA 96.37 372.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 372.455 97.14 372.825 ;
      VIA 96.37 372.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 372.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 367.035 97.16 367.365 ;
      VIA 96.37 367.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 367.015 97.14 367.385 ;
      VIA 96.37 367.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 367.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 361.595 97.16 361.925 ;
      VIA 96.37 361.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 361.575 97.14 361.945 ;
      VIA 96.37 361.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 361.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 356.155 97.16 356.485 ;
      VIA 96.37 356.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 356.135 97.14 356.505 ;
      VIA 96.37 356.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 356.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 350.715 97.16 351.045 ;
      VIA 96.37 350.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 350.695 97.14 351.065 ;
      VIA 96.37 350.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 350.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 345.275 97.16 345.605 ;
      VIA 96.37 345.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 345.255 97.14 345.625 ;
      VIA 96.37 345.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 345.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 339.835 97.16 340.165 ;
      VIA 96.37 340 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 339.815 97.14 340.185 ;
      VIA 96.37 340 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 340 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 334.395 97.16 334.725 ;
      VIA 96.37 334.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 334.375 97.14 334.745 ;
      VIA 96.37 334.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 334.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 328.955 97.16 329.285 ;
      VIA 96.37 329.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 328.935 97.14 329.305 ;
      VIA 96.37 329.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 329.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 323.515 97.16 323.845 ;
      VIA 96.37 323.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 323.495 97.14 323.865 ;
      VIA 96.37 323.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 323.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 318.075 97.16 318.405 ;
      VIA 96.37 318.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 318.055 97.14 318.425 ;
      VIA 96.37 318.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 318.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 312.635 97.16 312.965 ;
      VIA 96.37 312.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 312.615 97.14 312.985 ;
      VIA 96.37 312.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 312.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 307.195 97.16 307.525 ;
      VIA 96.37 307.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 307.175 97.14 307.545 ;
      VIA 96.37 307.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 307.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 301.755 97.16 302.085 ;
      VIA 96.37 301.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 301.735 97.14 302.105 ;
      VIA 96.37 301.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 301.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 296.315 97.16 296.645 ;
      VIA 96.37 296.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 296.295 97.14 296.665 ;
      VIA 96.37 296.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 296.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 290.875 97.16 291.205 ;
      VIA 96.37 291.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 290.855 97.14 291.225 ;
      VIA 96.37 291.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 291.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 285.435 97.16 285.765 ;
      VIA 96.37 285.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 285.415 97.14 285.785 ;
      VIA 96.37 285.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 285.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 279.995 97.16 280.325 ;
      VIA 96.37 280.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 279.975 97.14 280.345 ;
      VIA 96.37 280.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 280.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 274.555 97.16 274.885 ;
      VIA 96.37 274.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 274.535 97.14 274.905 ;
      VIA 96.37 274.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 274.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 269.115 97.16 269.445 ;
      VIA 96.37 269.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 269.095 97.14 269.465 ;
      VIA 96.37 269.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 269.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 263.675 97.16 264.005 ;
      VIA 96.37 263.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 263.655 97.14 264.025 ;
      VIA 96.37 263.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 263.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 258.235 97.16 258.565 ;
      VIA 96.37 258.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 258.215 97.14 258.585 ;
      VIA 96.37 258.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 258.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 252.795 97.16 253.125 ;
      VIA 96.37 252.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 252.775 97.14 253.145 ;
      VIA 96.37 252.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 252.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 247.355 97.16 247.685 ;
      VIA 96.37 247.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 247.335 97.14 247.705 ;
      VIA 96.37 247.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 247.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 241.915 97.16 242.245 ;
      VIA 96.37 242.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 241.895 97.14 242.265 ;
      VIA 96.37 242.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 242.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 236.475 97.16 236.805 ;
      VIA 96.37 236.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 236.455 97.14 236.825 ;
      VIA 96.37 236.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 236.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 231.035 97.16 231.365 ;
      VIA 96.37 231.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 231.015 97.14 231.385 ;
      VIA 96.37 231.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 231.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 225.595 97.16 225.925 ;
      VIA 96.37 225.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 225.575 97.14 225.945 ;
      VIA 96.37 225.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 225.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 220.155 97.16 220.485 ;
      VIA 96.37 220.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 220.135 97.14 220.505 ;
      VIA 96.37 220.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 220.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 214.715 97.16 215.045 ;
      VIA 96.37 214.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 214.695 97.14 215.065 ;
      VIA 96.37 214.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 214.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 209.275 97.16 209.605 ;
      VIA 96.37 209.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 209.255 97.14 209.625 ;
      VIA 96.37 209.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 209.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 203.835 97.16 204.165 ;
      VIA 96.37 204 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 203.815 97.14 204.185 ;
      VIA 96.37 204 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 204 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 198.395 97.16 198.725 ;
      VIA 96.37 198.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 198.375 97.14 198.745 ;
      VIA 96.37 198.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 198.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 192.955 97.16 193.285 ;
      VIA 96.37 193.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 192.935 97.14 193.305 ;
      VIA 96.37 193.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 193.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 187.515 97.16 187.845 ;
      VIA 96.37 187.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 187.495 97.14 187.865 ;
      VIA 96.37 187.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 187.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 182.075 97.16 182.405 ;
      VIA 96.37 182.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 182.055 97.14 182.425 ;
      VIA 96.37 182.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 182.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 176.635 97.16 176.965 ;
      VIA 96.37 176.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 176.615 97.14 176.985 ;
      VIA 96.37 176.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 176.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 171.195 97.16 171.525 ;
      VIA 96.37 171.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 171.175 97.14 171.545 ;
      VIA 96.37 171.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 171.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 165.755 97.16 166.085 ;
      VIA 96.37 165.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 165.735 97.14 166.105 ;
      VIA 96.37 165.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 165.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 160.315 97.16 160.645 ;
      VIA 96.37 160.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 160.295 97.14 160.665 ;
      VIA 96.37 160.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 160.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 154.875 97.16 155.205 ;
      VIA 96.37 155.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 154.855 97.14 155.225 ;
      VIA 96.37 155.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 155.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 149.435 97.16 149.765 ;
      VIA 96.37 149.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 149.415 97.14 149.785 ;
      VIA 96.37 149.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 149.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 143.995 97.16 144.325 ;
      VIA 96.37 144.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 143.975 97.14 144.345 ;
      VIA 96.37 144.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 144.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 138.555 97.16 138.885 ;
      VIA 96.37 138.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 138.535 97.14 138.905 ;
      VIA 96.37 138.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 138.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 133.115 97.16 133.445 ;
      VIA 96.37 133.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 133.095 97.14 133.465 ;
      VIA 96.37 133.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 133.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 127.675 97.16 128.005 ;
      VIA 96.37 127.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 127.655 97.14 128.025 ;
      VIA 96.37 127.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 127.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 122.235 97.16 122.565 ;
      VIA 96.37 122.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 122.215 97.14 122.585 ;
      VIA 96.37 122.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 122.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 116.795 97.16 117.125 ;
      VIA 96.37 116.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 116.775 97.14 117.145 ;
      VIA 96.37 116.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 116.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 111.355 97.16 111.685 ;
      VIA 96.37 111.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 111.335 97.14 111.705 ;
      VIA 96.37 111.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 111.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 105.915 97.16 106.245 ;
      VIA 96.37 106.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 105.895 97.14 106.265 ;
      VIA 96.37 106.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 106.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 100.475 97.16 100.805 ;
      VIA 96.37 100.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 100.455 97.14 100.825 ;
      VIA 96.37 100.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 100.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 95.035 97.16 95.365 ;
      VIA 96.37 95.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 95.015 97.14 95.385 ;
      VIA 96.37 95.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 95.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 89.595 97.16 89.925 ;
      VIA 96.37 89.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 89.575 97.14 89.945 ;
      VIA 96.37 89.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 89.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 84.155 97.16 84.485 ;
      VIA 96.37 84.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 84.135 97.14 84.505 ;
      VIA 96.37 84.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 84.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 78.715 97.16 79.045 ;
      VIA 96.37 78.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 78.695 97.14 79.065 ;
      VIA 96.37 78.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 78.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 73.275 97.16 73.605 ;
      VIA 96.37 73.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 73.255 97.14 73.625 ;
      VIA 96.37 73.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 73.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 67.835 97.16 68.165 ;
      VIA 96.37 68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 67.815 97.14 68.185 ;
      VIA 96.37 68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 62.395 97.16 62.725 ;
      VIA 96.37 62.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 62.375 97.14 62.745 ;
      VIA 96.37 62.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 62.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 56.955 97.16 57.285 ;
      VIA 96.37 57.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 56.935 97.14 57.305 ;
      VIA 96.37 57.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 57.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 51.515 97.16 51.845 ;
      VIA 96.37 51.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 51.495 97.14 51.865 ;
      VIA 96.37 51.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 51.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 46.075 97.16 46.405 ;
      VIA 96.37 46.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 46.055 97.14 46.425 ;
      VIA 96.37 46.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 46.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 40.635 97.16 40.965 ;
      VIA 96.37 40.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 40.615 97.14 40.985 ;
      VIA 96.37 40.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 40.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 35.195 97.16 35.525 ;
      VIA 96.37 35.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 35.175 97.14 35.545 ;
      VIA 96.37 35.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 35.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 29.755 97.16 30.085 ;
      VIA 96.37 29.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 29.735 97.14 30.105 ;
      VIA 96.37 29.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 29.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 24.315 97.16 24.645 ;
      VIA 96.37 24.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 24.295 97.14 24.665 ;
      VIA 96.37 24.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 24.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 18.875 97.16 19.205 ;
      VIA 96.37 19.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 18.855 97.14 19.225 ;
      VIA 96.37 19.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 19.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 13.435 97.16 13.765 ;
      VIA 96.37 13.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 13.415 97.14 13.785 ;
      VIA 96.37 13.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 13.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 7.995 97.16 8.325 ;
      VIA 96.37 8.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 7.975 97.14 8.345 ;
      VIA 96.37 8.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 8.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  95.58 2.555 97.16 2.885 ;
      VIA 96.37 2.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  95.6 2.535 97.14 2.905 ;
      VIA 96.37 2.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 96.37 2.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 698.875 70.02 699.205 ;
      VIA 69.23 699.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 698.855 70 699.225 ;
      VIA 69.23 699.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 699.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 693.435 70.02 693.765 ;
      VIA 69.23 693.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 693.415 70 693.785 ;
      VIA 69.23 693.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 693.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 687.995 70.02 688.325 ;
      VIA 69.23 688.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 687.975 70 688.345 ;
      VIA 69.23 688.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 688.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 682.555 70.02 682.885 ;
      VIA 69.23 682.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 682.535 70 682.905 ;
      VIA 69.23 682.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 682.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 677.115 70.02 677.445 ;
      VIA 69.23 677.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 677.095 70 677.465 ;
      VIA 69.23 677.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 677.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 671.675 70.02 672.005 ;
      VIA 69.23 671.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 671.655 70 672.025 ;
      VIA 69.23 671.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 671.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 666.235 70.02 666.565 ;
      VIA 69.23 666.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 666.215 70 666.585 ;
      VIA 69.23 666.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 666.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 660.795 70.02 661.125 ;
      VIA 69.23 660.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 660.775 70 661.145 ;
      VIA 69.23 660.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 660.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 655.355 70.02 655.685 ;
      VIA 69.23 655.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 655.335 70 655.705 ;
      VIA 69.23 655.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 655.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 649.915 70.02 650.245 ;
      VIA 69.23 650.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 649.895 70 650.265 ;
      VIA 69.23 650.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 650.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 644.475 70.02 644.805 ;
      VIA 69.23 644.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 644.455 70 644.825 ;
      VIA 69.23 644.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 644.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 639.035 70.02 639.365 ;
      VIA 69.23 639.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 639.015 70 639.385 ;
      VIA 69.23 639.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 639.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 633.595 70.02 633.925 ;
      VIA 69.23 633.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 633.575 70 633.945 ;
      VIA 69.23 633.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 633.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 628.155 70.02 628.485 ;
      VIA 69.23 628.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 628.135 70 628.505 ;
      VIA 69.23 628.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 628.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 622.715 70.02 623.045 ;
      VIA 69.23 622.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 622.695 70 623.065 ;
      VIA 69.23 622.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 622.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 617.275 70.02 617.605 ;
      VIA 69.23 617.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 617.255 70 617.625 ;
      VIA 69.23 617.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 617.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 611.835 70.02 612.165 ;
      VIA 69.23 612 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 611.815 70 612.185 ;
      VIA 69.23 612 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 612 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 606.395 70.02 606.725 ;
      VIA 69.23 606.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 606.375 70 606.745 ;
      VIA 69.23 606.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 606.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 600.955 70.02 601.285 ;
      VIA 69.23 601.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 600.935 70 601.305 ;
      VIA 69.23 601.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 601.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 595.515 70.02 595.845 ;
      VIA 69.23 595.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 595.495 70 595.865 ;
      VIA 69.23 595.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 595.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 590.075 70.02 590.405 ;
      VIA 69.23 590.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 590.055 70 590.425 ;
      VIA 69.23 590.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 590.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 584.635 70.02 584.965 ;
      VIA 69.23 584.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 584.615 70 584.985 ;
      VIA 69.23 584.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 584.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 579.195 70.02 579.525 ;
      VIA 69.23 579.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 579.175 70 579.545 ;
      VIA 69.23 579.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 579.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 573.755 70.02 574.085 ;
      VIA 69.23 573.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 573.735 70 574.105 ;
      VIA 69.23 573.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 573.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 568.315 70.02 568.645 ;
      VIA 69.23 568.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 568.295 70 568.665 ;
      VIA 69.23 568.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 568.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 562.875 70.02 563.205 ;
      VIA 69.23 563.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 562.855 70 563.225 ;
      VIA 69.23 563.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 563.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 557.435 70.02 557.765 ;
      VIA 69.23 557.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 557.415 70 557.785 ;
      VIA 69.23 557.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 557.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 551.995 70.02 552.325 ;
      VIA 69.23 552.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 551.975 70 552.345 ;
      VIA 69.23 552.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 552.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 546.555 70.02 546.885 ;
      VIA 69.23 546.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 546.535 70 546.905 ;
      VIA 69.23 546.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 546.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 541.115 70.02 541.445 ;
      VIA 69.23 541.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 541.095 70 541.465 ;
      VIA 69.23 541.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 541.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 535.675 70.02 536.005 ;
      VIA 69.23 535.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 535.655 70 536.025 ;
      VIA 69.23 535.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 535.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 530.235 70.02 530.565 ;
      VIA 69.23 530.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 530.215 70 530.585 ;
      VIA 69.23 530.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 530.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 524.795 70.02 525.125 ;
      VIA 69.23 524.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 524.775 70 525.145 ;
      VIA 69.23 524.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 524.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 519.355 70.02 519.685 ;
      VIA 69.23 519.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 519.335 70 519.705 ;
      VIA 69.23 519.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 519.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 513.915 70.02 514.245 ;
      VIA 69.23 514.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 513.895 70 514.265 ;
      VIA 69.23 514.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 514.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 508.475 70.02 508.805 ;
      VIA 69.23 508.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 508.455 70 508.825 ;
      VIA 69.23 508.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 508.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 503.035 70.02 503.365 ;
      VIA 69.23 503.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 503.015 70 503.385 ;
      VIA 69.23 503.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 503.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 497.595 70.02 497.925 ;
      VIA 69.23 497.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 497.575 70 497.945 ;
      VIA 69.23 497.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 497.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 492.155 70.02 492.485 ;
      VIA 69.23 492.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 492.135 70 492.505 ;
      VIA 69.23 492.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 492.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 486.715 70.02 487.045 ;
      VIA 69.23 486.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 486.695 70 487.065 ;
      VIA 69.23 486.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 486.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 481.275 70.02 481.605 ;
      VIA 69.23 481.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 481.255 70 481.625 ;
      VIA 69.23 481.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 481.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 475.835 70.02 476.165 ;
      VIA 69.23 476 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 475.815 70 476.185 ;
      VIA 69.23 476 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 476 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 470.395 70.02 470.725 ;
      VIA 69.23 470.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 470.375 70 470.745 ;
      VIA 69.23 470.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 470.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 464.955 70.02 465.285 ;
      VIA 69.23 465.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 464.935 70 465.305 ;
      VIA 69.23 465.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 465.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 459.515 70.02 459.845 ;
      VIA 69.23 459.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 459.495 70 459.865 ;
      VIA 69.23 459.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 459.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 454.075 70.02 454.405 ;
      VIA 69.23 454.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 454.055 70 454.425 ;
      VIA 69.23 454.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 454.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 448.635 70.02 448.965 ;
      VIA 69.23 448.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 448.615 70 448.985 ;
      VIA 69.23 448.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 448.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 443.195 70.02 443.525 ;
      VIA 69.23 443.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 443.175 70 443.545 ;
      VIA 69.23 443.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 443.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 437.755 70.02 438.085 ;
      VIA 69.23 437.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 437.735 70 438.105 ;
      VIA 69.23 437.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 437.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 432.315 70.02 432.645 ;
      VIA 69.23 432.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 432.295 70 432.665 ;
      VIA 69.23 432.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 432.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 426.875 70.02 427.205 ;
      VIA 69.23 427.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 426.855 70 427.225 ;
      VIA 69.23 427.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 427.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 421.435 70.02 421.765 ;
      VIA 69.23 421.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 421.415 70 421.785 ;
      VIA 69.23 421.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 421.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 415.995 70.02 416.325 ;
      VIA 69.23 416.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 415.975 70 416.345 ;
      VIA 69.23 416.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 416.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 410.555 70.02 410.885 ;
      VIA 69.23 410.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 410.535 70 410.905 ;
      VIA 69.23 410.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 410.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 405.115 70.02 405.445 ;
      VIA 69.23 405.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 405.095 70 405.465 ;
      VIA 69.23 405.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 405.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 399.675 70.02 400.005 ;
      VIA 69.23 399.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 399.655 70 400.025 ;
      VIA 69.23 399.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 399.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 394.235 70.02 394.565 ;
      VIA 69.23 394.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 394.215 70 394.585 ;
      VIA 69.23 394.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 394.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 388.795 70.02 389.125 ;
      VIA 69.23 388.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 388.775 70 389.145 ;
      VIA 69.23 388.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 388.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 383.355 70.02 383.685 ;
      VIA 69.23 383.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 383.335 70 383.705 ;
      VIA 69.23 383.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 383.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 377.915 70.02 378.245 ;
      VIA 69.23 378.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 377.895 70 378.265 ;
      VIA 69.23 378.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 378.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 372.475 70.02 372.805 ;
      VIA 69.23 372.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 372.455 70 372.825 ;
      VIA 69.23 372.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 372.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 367.035 70.02 367.365 ;
      VIA 69.23 367.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 367.015 70 367.385 ;
      VIA 69.23 367.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 367.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 361.595 70.02 361.925 ;
      VIA 69.23 361.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 361.575 70 361.945 ;
      VIA 69.23 361.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 361.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 356.155 70.02 356.485 ;
      VIA 69.23 356.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 356.135 70 356.505 ;
      VIA 69.23 356.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 356.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 350.715 70.02 351.045 ;
      VIA 69.23 350.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 350.695 70 351.065 ;
      VIA 69.23 350.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 350.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 345.275 70.02 345.605 ;
      VIA 69.23 345.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 345.255 70 345.625 ;
      VIA 69.23 345.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 345.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 339.835 70.02 340.165 ;
      VIA 69.23 340 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 339.815 70 340.185 ;
      VIA 69.23 340 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 340 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 334.395 70.02 334.725 ;
      VIA 69.23 334.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 334.375 70 334.745 ;
      VIA 69.23 334.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 334.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 328.955 70.02 329.285 ;
      VIA 69.23 329.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 328.935 70 329.305 ;
      VIA 69.23 329.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 329.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 323.515 70.02 323.845 ;
      VIA 69.23 323.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 323.495 70 323.865 ;
      VIA 69.23 323.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 323.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 318.075 70.02 318.405 ;
      VIA 69.23 318.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 318.055 70 318.425 ;
      VIA 69.23 318.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 318.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 312.635 70.02 312.965 ;
      VIA 69.23 312.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 312.615 70 312.985 ;
      VIA 69.23 312.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 312.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 307.195 70.02 307.525 ;
      VIA 69.23 307.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 307.175 70 307.545 ;
      VIA 69.23 307.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 307.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 301.755 70.02 302.085 ;
      VIA 69.23 301.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 301.735 70 302.105 ;
      VIA 69.23 301.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 301.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 296.315 70.02 296.645 ;
      VIA 69.23 296.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 296.295 70 296.665 ;
      VIA 69.23 296.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 296.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 290.875 70.02 291.205 ;
      VIA 69.23 291.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 290.855 70 291.225 ;
      VIA 69.23 291.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 291.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 285.435 70.02 285.765 ;
      VIA 69.23 285.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 285.415 70 285.785 ;
      VIA 69.23 285.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 285.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 279.995 70.02 280.325 ;
      VIA 69.23 280.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 279.975 70 280.345 ;
      VIA 69.23 280.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 280.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 274.555 70.02 274.885 ;
      VIA 69.23 274.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 274.535 70 274.905 ;
      VIA 69.23 274.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 274.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 269.115 70.02 269.445 ;
      VIA 69.23 269.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 269.095 70 269.465 ;
      VIA 69.23 269.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 269.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 263.675 70.02 264.005 ;
      VIA 69.23 263.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 263.655 70 264.025 ;
      VIA 69.23 263.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 263.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 258.235 70.02 258.565 ;
      VIA 69.23 258.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 258.215 70 258.585 ;
      VIA 69.23 258.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 258.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 252.795 70.02 253.125 ;
      VIA 69.23 252.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 252.775 70 253.145 ;
      VIA 69.23 252.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 252.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 247.355 70.02 247.685 ;
      VIA 69.23 247.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 247.335 70 247.705 ;
      VIA 69.23 247.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 247.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 241.915 70.02 242.245 ;
      VIA 69.23 242.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 241.895 70 242.265 ;
      VIA 69.23 242.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 242.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 236.475 70.02 236.805 ;
      VIA 69.23 236.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 236.455 70 236.825 ;
      VIA 69.23 236.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 236.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 231.035 70.02 231.365 ;
      VIA 69.23 231.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 231.015 70 231.385 ;
      VIA 69.23 231.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 231.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 225.595 70.02 225.925 ;
      VIA 69.23 225.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 225.575 70 225.945 ;
      VIA 69.23 225.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 225.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 220.155 70.02 220.485 ;
      VIA 69.23 220.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 220.135 70 220.505 ;
      VIA 69.23 220.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 220.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 214.715 70.02 215.045 ;
      VIA 69.23 214.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 214.695 70 215.065 ;
      VIA 69.23 214.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 214.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 209.275 70.02 209.605 ;
      VIA 69.23 209.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 209.255 70 209.625 ;
      VIA 69.23 209.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 209.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 203.835 70.02 204.165 ;
      VIA 69.23 204 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 203.815 70 204.185 ;
      VIA 69.23 204 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 204 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 198.395 70.02 198.725 ;
      VIA 69.23 198.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 198.375 70 198.745 ;
      VIA 69.23 198.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 198.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 192.955 70.02 193.285 ;
      VIA 69.23 193.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 192.935 70 193.305 ;
      VIA 69.23 193.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 193.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 187.515 70.02 187.845 ;
      VIA 69.23 187.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 187.495 70 187.865 ;
      VIA 69.23 187.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 187.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 182.075 70.02 182.405 ;
      VIA 69.23 182.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 182.055 70 182.425 ;
      VIA 69.23 182.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 182.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 176.635 70.02 176.965 ;
      VIA 69.23 176.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 176.615 70 176.985 ;
      VIA 69.23 176.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 176.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 171.195 70.02 171.525 ;
      VIA 69.23 171.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 171.175 70 171.545 ;
      VIA 69.23 171.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 171.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 165.755 70.02 166.085 ;
      VIA 69.23 165.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 165.735 70 166.105 ;
      VIA 69.23 165.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 165.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 160.315 70.02 160.645 ;
      VIA 69.23 160.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 160.295 70 160.665 ;
      VIA 69.23 160.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 160.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 154.875 70.02 155.205 ;
      VIA 69.23 155.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 154.855 70 155.225 ;
      VIA 69.23 155.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 155.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 149.435 70.02 149.765 ;
      VIA 69.23 149.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 149.415 70 149.785 ;
      VIA 69.23 149.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 149.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 143.995 70.02 144.325 ;
      VIA 69.23 144.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 143.975 70 144.345 ;
      VIA 69.23 144.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 144.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 138.555 70.02 138.885 ;
      VIA 69.23 138.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 138.535 70 138.905 ;
      VIA 69.23 138.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 138.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 133.115 70.02 133.445 ;
      VIA 69.23 133.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 133.095 70 133.465 ;
      VIA 69.23 133.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 133.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 127.675 70.02 128.005 ;
      VIA 69.23 127.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 127.655 70 128.025 ;
      VIA 69.23 127.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 127.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 122.235 70.02 122.565 ;
      VIA 69.23 122.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 122.215 70 122.585 ;
      VIA 69.23 122.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 122.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 116.795 70.02 117.125 ;
      VIA 69.23 116.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 116.775 70 117.145 ;
      VIA 69.23 116.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 116.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 111.355 70.02 111.685 ;
      VIA 69.23 111.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 111.335 70 111.705 ;
      VIA 69.23 111.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 111.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 105.915 70.02 106.245 ;
      VIA 69.23 106.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 105.895 70 106.265 ;
      VIA 69.23 106.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 106.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 100.475 70.02 100.805 ;
      VIA 69.23 100.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 100.455 70 100.825 ;
      VIA 69.23 100.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 100.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 95.035 70.02 95.365 ;
      VIA 69.23 95.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 95.015 70 95.385 ;
      VIA 69.23 95.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 95.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 89.595 70.02 89.925 ;
      VIA 69.23 89.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 89.575 70 89.945 ;
      VIA 69.23 89.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 89.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 84.155 70.02 84.485 ;
      VIA 69.23 84.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 84.135 70 84.505 ;
      VIA 69.23 84.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 84.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 78.715 70.02 79.045 ;
      VIA 69.23 78.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 78.695 70 79.065 ;
      VIA 69.23 78.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 78.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 73.275 70.02 73.605 ;
      VIA 69.23 73.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 73.255 70 73.625 ;
      VIA 69.23 73.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 73.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 67.835 70.02 68.165 ;
      VIA 69.23 68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 67.815 70 68.185 ;
      VIA 69.23 68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 62.395 70.02 62.725 ;
      VIA 69.23 62.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 62.375 70 62.745 ;
      VIA 69.23 62.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 62.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 56.955 70.02 57.285 ;
      VIA 69.23 57.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 56.935 70 57.305 ;
      VIA 69.23 57.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 57.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 51.515 70.02 51.845 ;
      VIA 69.23 51.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 51.495 70 51.865 ;
      VIA 69.23 51.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 51.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 46.075 70.02 46.405 ;
      VIA 69.23 46.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 46.055 70 46.425 ;
      VIA 69.23 46.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 46.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 40.635 70.02 40.965 ;
      VIA 69.23 40.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 40.615 70 40.985 ;
      VIA 69.23 40.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 40.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 35.195 70.02 35.525 ;
      VIA 69.23 35.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 35.175 70 35.545 ;
      VIA 69.23 35.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 35.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 29.755 70.02 30.085 ;
      VIA 69.23 29.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 29.735 70 30.105 ;
      VIA 69.23 29.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 29.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 24.315 70.02 24.645 ;
      VIA 69.23 24.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 24.295 70 24.665 ;
      VIA 69.23 24.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 24.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 18.875 70.02 19.205 ;
      VIA 69.23 19.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 18.855 70 19.225 ;
      VIA 69.23 19.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 19.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 13.435 70.02 13.765 ;
      VIA 69.23 13.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 13.415 70 13.785 ;
      VIA 69.23 13.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 13.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 7.995 70.02 8.325 ;
      VIA 69.23 8.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 7.975 70 8.345 ;
      VIA 69.23 8.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 8.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  68.44 2.555 70.02 2.885 ;
      VIA 69.23 2.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  68.46 2.535 70 2.905 ;
      VIA 69.23 2.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 69.23 2.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 698.875 42.88 699.205 ;
      VIA 42.09 699.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 698.855 42.86 699.225 ;
      VIA 42.09 699.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 699.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 693.435 42.88 693.765 ;
      VIA 42.09 693.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 693.415 42.86 693.785 ;
      VIA 42.09 693.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 693.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 687.995 42.88 688.325 ;
      VIA 42.09 688.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 687.975 42.86 688.345 ;
      VIA 42.09 688.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 688.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 682.555 42.88 682.885 ;
      VIA 42.09 682.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 682.535 42.86 682.905 ;
      VIA 42.09 682.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 682.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 677.115 42.88 677.445 ;
      VIA 42.09 677.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 677.095 42.86 677.465 ;
      VIA 42.09 677.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 677.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 671.675 42.88 672.005 ;
      VIA 42.09 671.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 671.655 42.86 672.025 ;
      VIA 42.09 671.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 671.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 666.235 42.88 666.565 ;
      VIA 42.09 666.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 666.215 42.86 666.585 ;
      VIA 42.09 666.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 666.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 660.795 42.88 661.125 ;
      VIA 42.09 660.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 660.775 42.86 661.145 ;
      VIA 42.09 660.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 660.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 655.355 42.88 655.685 ;
      VIA 42.09 655.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 655.335 42.86 655.705 ;
      VIA 42.09 655.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 655.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 649.915 42.88 650.245 ;
      VIA 42.09 650.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 649.895 42.86 650.265 ;
      VIA 42.09 650.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 650.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 644.475 42.88 644.805 ;
      VIA 42.09 644.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 644.455 42.86 644.825 ;
      VIA 42.09 644.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 644.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 639.035 42.88 639.365 ;
      VIA 42.09 639.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 639.015 42.86 639.385 ;
      VIA 42.09 639.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 639.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 633.595 42.88 633.925 ;
      VIA 42.09 633.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 633.575 42.86 633.945 ;
      VIA 42.09 633.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 633.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 628.155 42.88 628.485 ;
      VIA 42.09 628.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 628.135 42.86 628.505 ;
      VIA 42.09 628.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 628.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 622.715 42.88 623.045 ;
      VIA 42.09 622.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 622.695 42.86 623.065 ;
      VIA 42.09 622.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 622.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 617.275 42.88 617.605 ;
      VIA 42.09 617.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 617.255 42.86 617.625 ;
      VIA 42.09 617.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 617.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 611.835 42.88 612.165 ;
      VIA 42.09 612 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 611.815 42.86 612.185 ;
      VIA 42.09 612 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 612 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 606.395 42.88 606.725 ;
      VIA 42.09 606.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 606.375 42.86 606.745 ;
      VIA 42.09 606.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 606.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 600.955 42.88 601.285 ;
      VIA 42.09 601.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 600.935 42.86 601.305 ;
      VIA 42.09 601.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 601.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 595.515 42.88 595.845 ;
      VIA 42.09 595.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 595.495 42.86 595.865 ;
      VIA 42.09 595.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 595.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 590.075 42.88 590.405 ;
      VIA 42.09 590.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 590.055 42.86 590.425 ;
      VIA 42.09 590.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 590.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 584.635 42.88 584.965 ;
      VIA 42.09 584.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 584.615 42.86 584.985 ;
      VIA 42.09 584.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 584.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 579.195 42.88 579.525 ;
      VIA 42.09 579.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 579.175 42.86 579.545 ;
      VIA 42.09 579.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 579.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 573.755 42.88 574.085 ;
      VIA 42.09 573.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 573.735 42.86 574.105 ;
      VIA 42.09 573.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 573.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 568.315 42.88 568.645 ;
      VIA 42.09 568.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 568.295 42.86 568.665 ;
      VIA 42.09 568.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 568.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 562.875 42.88 563.205 ;
      VIA 42.09 563.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 562.855 42.86 563.225 ;
      VIA 42.09 563.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 563.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 557.435 42.88 557.765 ;
      VIA 42.09 557.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 557.415 42.86 557.785 ;
      VIA 42.09 557.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 557.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 551.995 42.88 552.325 ;
      VIA 42.09 552.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 551.975 42.86 552.345 ;
      VIA 42.09 552.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 552.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 546.555 42.88 546.885 ;
      VIA 42.09 546.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 546.535 42.86 546.905 ;
      VIA 42.09 546.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 546.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 541.115 42.88 541.445 ;
      VIA 42.09 541.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 541.095 42.86 541.465 ;
      VIA 42.09 541.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 541.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 535.675 42.88 536.005 ;
      VIA 42.09 535.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 535.655 42.86 536.025 ;
      VIA 42.09 535.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 535.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 530.235 42.88 530.565 ;
      VIA 42.09 530.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 530.215 42.86 530.585 ;
      VIA 42.09 530.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 530.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 524.795 42.88 525.125 ;
      VIA 42.09 524.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 524.775 42.86 525.145 ;
      VIA 42.09 524.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 524.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 519.355 42.88 519.685 ;
      VIA 42.09 519.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 519.335 42.86 519.705 ;
      VIA 42.09 519.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 519.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 513.915 42.88 514.245 ;
      VIA 42.09 514.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 513.895 42.86 514.265 ;
      VIA 42.09 514.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 514.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 508.475 42.88 508.805 ;
      VIA 42.09 508.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 508.455 42.86 508.825 ;
      VIA 42.09 508.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 508.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 503.035 42.88 503.365 ;
      VIA 42.09 503.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 503.015 42.86 503.385 ;
      VIA 42.09 503.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 503.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 497.595 42.88 497.925 ;
      VIA 42.09 497.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 497.575 42.86 497.945 ;
      VIA 42.09 497.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 497.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 492.155 42.88 492.485 ;
      VIA 42.09 492.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 492.135 42.86 492.505 ;
      VIA 42.09 492.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 492.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 486.715 42.88 487.045 ;
      VIA 42.09 486.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 486.695 42.86 487.065 ;
      VIA 42.09 486.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 486.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 481.275 42.88 481.605 ;
      VIA 42.09 481.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 481.255 42.86 481.625 ;
      VIA 42.09 481.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 481.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 475.835 42.88 476.165 ;
      VIA 42.09 476 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 475.815 42.86 476.185 ;
      VIA 42.09 476 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 476 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 470.395 42.88 470.725 ;
      VIA 42.09 470.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 470.375 42.86 470.745 ;
      VIA 42.09 470.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 470.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 464.955 42.88 465.285 ;
      VIA 42.09 465.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 464.935 42.86 465.305 ;
      VIA 42.09 465.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 465.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 459.515 42.88 459.845 ;
      VIA 42.09 459.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 459.495 42.86 459.865 ;
      VIA 42.09 459.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 459.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 454.075 42.88 454.405 ;
      VIA 42.09 454.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 454.055 42.86 454.425 ;
      VIA 42.09 454.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 454.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 448.635 42.88 448.965 ;
      VIA 42.09 448.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 448.615 42.86 448.985 ;
      VIA 42.09 448.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 448.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 443.195 42.88 443.525 ;
      VIA 42.09 443.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 443.175 42.86 443.545 ;
      VIA 42.09 443.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 443.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 437.755 42.88 438.085 ;
      VIA 42.09 437.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 437.735 42.86 438.105 ;
      VIA 42.09 437.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 437.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 432.315 42.88 432.645 ;
      VIA 42.09 432.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 432.295 42.86 432.665 ;
      VIA 42.09 432.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 432.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 426.875 42.88 427.205 ;
      VIA 42.09 427.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 426.855 42.86 427.225 ;
      VIA 42.09 427.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 427.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 421.435 42.88 421.765 ;
      VIA 42.09 421.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 421.415 42.86 421.785 ;
      VIA 42.09 421.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 421.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 415.995 42.88 416.325 ;
      VIA 42.09 416.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 415.975 42.86 416.345 ;
      VIA 42.09 416.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 416.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 410.555 42.88 410.885 ;
      VIA 42.09 410.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 410.535 42.86 410.905 ;
      VIA 42.09 410.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 410.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 405.115 42.88 405.445 ;
      VIA 42.09 405.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 405.095 42.86 405.465 ;
      VIA 42.09 405.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 405.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 399.675 42.88 400.005 ;
      VIA 42.09 399.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 399.655 42.86 400.025 ;
      VIA 42.09 399.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 399.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 394.235 42.88 394.565 ;
      VIA 42.09 394.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 394.215 42.86 394.585 ;
      VIA 42.09 394.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 394.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 388.795 42.88 389.125 ;
      VIA 42.09 388.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 388.775 42.86 389.145 ;
      VIA 42.09 388.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 388.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 383.355 42.88 383.685 ;
      VIA 42.09 383.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 383.335 42.86 383.705 ;
      VIA 42.09 383.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 383.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 377.915 42.88 378.245 ;
      VIA 42.09 378.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 377.895 42.86 378.265 ;
      VIA 42.09 378.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 378.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 372.475 42.88 372.805 ;
      VIA 42.09 372.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 372.455 42.86 372.825 ;
      VIA 42.09 372.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 372.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 367.035 42.88 367.365 ;
      VIA 42.09 367.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 367.015 42.86 367.385 ;
      VIA 42.09 367.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 367.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 361.595 42.88 361.925 ;
      VIA 42.09 361.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 361.575 42.86 361.945 ;
      VIA 42.09 361.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 361.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 356.155 42.88 356.485 ;
      VIA 42.09 356.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 356.135 42.86 356.505 ;
      VIA 42.09 356.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 356.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 350.715 42.88 351.045 ;
      VIA 42.09 350.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 350.695 42.86 351.065 ;
      VIA 42.09 350.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 350.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 345.275 42.88 345.605 ;
      VIA 42.09 345.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 345.255 42.86 345.625 ;
      VIA 42.09 345.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 345.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 339.835 42.88 340.165 ;
      VIA 42.09 340 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 339.815 42.86 340.185 ;
      VIA 42.09 340 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 340 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 334.395 42.88 334.725 ;
      VIA 42.09 334.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 334.375 42.86 334.745 ;
      VIA 42.09 334.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 334.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 328.955 42.88 329.285 ;
      VIA 42.09 329.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 328.935 42.86 329.305 ;
      VIA 42.09 329.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 329.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 323.515 42.88 323.845 ;
      VIA 42.09 323.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 323.495 42.86 323.865 ;
      VIA 42.09 323.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 323.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 318.075 42.88 318.405 ;
      VIA 42.09 318.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 318.055 42.86 318.425 ;
      VIA 42.09 318.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 318.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 312.635 42.88 312.965 ;
      VIA 42.09 312.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 312.615 42.86 312.985 ;
      VIA 42.09 312.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 312.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 307.195 42.88 307.525 ;
      VIA 42.09 307.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 307.175 42.86 307.545 ;
      VIA 42.09 307.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 307.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 301.755 42.88 302.085 ;
      VIA 42.09 301.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 301.735 42.86 302.105 ;
      VIA 42.09 301.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 301.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 296.315 42.88 296.645 ;
      VIA 42.09 296.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 296.295 42.86 296.665 ;
      VIA 42.09 296.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 296.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 290.875 42.88 291.205 ;
      VIA 42.09 291.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 290.855 42.86 291.225 ;
      VIA 42.09 291.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 291.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 285.435 42.88 285.765 ;
      VIA 42.09 285.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 285.415 42.86 285.785 ;
      VIA 42.09 285.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 285.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 279.995 42.88 280.325 ;
      VIA 42.09 280.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 279.975 42.86 280.345 ;
      VIA 42.09 280.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 280.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 274.555 42.88 274.885 ;
      VIA 42.09 274.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 274.535 42.86 274.905 ;
      VIA 42.09 274.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 274.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 269.115 42.88 269.445 ;
      VIA 42.09 269.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 269.095 42.86 269.465 ;
      VIA 42.09 269.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 269.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 263.675 42.88 264.005 ;
      VIA 42.09 263.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 263.655 42.86 264.025 ;
      VIA 42.09 263.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 263.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 258.235 42.88 258.565 ;
      VIA 42.09 258.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 258.215 42.86 258.585 ;
      VIA 42.09 258.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 258.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 252.795 42.88 253.125 ;
      VIA 42.09 252.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 252.775 42.86 253.145 ;
      VIA 42.09 252.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 252.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 247.355 42.88 247.685 ;
      VIA 42.09 247.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 247.335 42.86 247.705 ;
      VIA 42.09 247.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 247.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 241.915 42.88 242.245 ;
      VIA 42.09 242.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 241.895 42.86 242.265 ;
      VIA 42.09 242.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 242.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 236.475 42.88 236.805 ;
      VIA 42.09 236.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 236.455 42.86 236.825 ;
      VIA 42.09 236.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 236.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 231.035 42.88 231.365 ;
      VIA 42.09 231.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 231.015 42.86 231.385 ;
      VIA 42.09 231.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 231.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 225.595 42.88 225.925 ;
      VIA 42.09 225.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 225.575 42.86 225.945 ;
      VIA 42.09 225.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 225.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 220.155 42.88 220.485 ;
      VIA 42.09 220.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 220.135 42.86 220.505 ;
      VIA 42.09 220.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 220.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 214.715 42.88 215.045 ;
      VIA 42.09 214.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 214.695 42.86 215.065 ;
      VIA 42.09 214.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 214.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 209.275 42.88 209.605 ;
      VIA 42.09 209.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 209.255 42.86 209.625 ;
      VIA 42.09 209.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 209.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 203.835 42.88 204.165 ;
      VIA 42.09 204 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 203.815 42.86 204.185 ;
      VIA 42.09 204 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 204 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 198.395 42.88 198.725 ;
      VIA 42.09 198.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 198.375 42.86 198.745 ;
      VIA 42.09 198.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 198.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 192.955 42.88 193.285 ;
      VIA 42.09 193.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 192.935 42.86 193.305 ;
      VIA 42.09 193.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 193.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 187.515 42.88 187.845 ;
      VIA 42.09 187.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 187.495 42.86 187.865 ;
      VIA 42.09 187.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 187.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 182.075 42.88 182.405 ;
      VIA 42.09 182.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 182.055 42.86 182.425 ;
      VIA 42.09 182.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 182.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 176.635 42.88 176.965 ;
      VIA 42.09 176.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 176.615 42.86 176.985 ;
      VIA 42.09 176.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 176.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 171.195 42.88 171.525 ;
      VIA 42.09 171.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 171.175 42.86 171.545 ;
      VIA 42.09 171.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 171.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 165.755 42.88 166.085 ;
      VIA 42.09 165.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 165.735 42.86 166.105 ;
      VIA 42.09 165.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 165.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 160.315 42.88 160.645 ;
      VIA 42.09 160.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 160.295 42.86 160.665 ;
      VIA 42.09 160.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 160.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 154.875 42.88 155.205 ;
      VIA 42.09 155.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 154.855 42.86 155.225 ;
      VIA 42.09 155.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 155.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 149.435 42.88 149.765 ;
      VIA 42.09 149.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 149.415 42.86 149.785 ;
      VIA 42.09 149.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 149.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 143.995 42.88 144.325 ;
      VIA 42.09 144.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 143.975 42.86 144.345 ;
      VIA 42.09 144.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 144.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 138.555 42.88 138.885 ;
      VIA 42.09 138.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 138.535 42.86 138.905 ;
      VIA 42.09 138.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 138.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 133.115 42.88 133.445 ;
      VIA 42.09 133.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 133.095 42.86 133.465 ;
      VIA 42.09 133.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 133.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 127.675 42.88 128.005 ;
      VIA 42.09 127.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 127.655 42.86 128.025 ;
      VIA 42.09 127.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 127.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 122.235 42.88 122.565 ;
      VIA 42.09 122.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 122.215 42.86 122.585 ;
      VIA 42.09 122.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 122.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 116.795 42.88 117.125 ;
      VIA 42.09 116.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 116.775 42.86 117.145 ;
      VIA 42.09 116.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 116.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 111.355 42.88 111.685 ;
      VIA 42.09 111.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 111.335 42.86 111.705 ;
      VIA 42.09 111.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 111.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 105.915 42.88 106.245 ;
      VIA 42.09 106.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 105.895 42.86 106.265 ;
      VIA 42.09 106.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 106.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 100.475 42.88 100.805 ;
      VIA 42.09 100.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 100.455 42.86 100.825 ;
      VIA 42.09 100.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 100.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 95.035 42.88 95.365 ;
      VIA 42.09 95.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 95.015 42.86 95.385 ;
      VIA 42.09 95.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 95.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 89.595 42.88 89.925 ;
      VIA 42.09 89.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 89.575 42.86 89.945 ;
      VIA 42.09 89.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 89.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 84.155 42.88 84.485 ;
      VIA 42.09 84.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 84.135 42.86 84.505 ;
      VIA 42.09 84.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 84.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 78.715 42.88 79.045 ;
      VIA 42.09 78.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 78.695 42.86 79.065 ;
      VIA 42.09 78.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 78.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 73.275 42.88 73.605 ;
      VIA 42.09 73.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 73.255 42.86 73.625 ;
      VIA 42.09 73.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 73.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 67.835 42.88 68.165 ;
      VIA 42.09 68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 67.815 42.86 68.185 ;
      VIA 42.09 68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 62.395 42.88 62.725 ;
      VIA 42.09 62.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 62.375 42.86 62.745 ;
      VIA 42.09 62.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 62.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 56.955 42.88 57.285 ;
      VIA 42.09 57.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 56.935 42.86 57.305 ;
      VIA 42.09 57.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 57.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 51.515 42.88 51.845 ;
      VIA 42.09 51.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 51.495 42.86 51.865 ;
      VIA 42.09 51.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 51.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 46.075 42.88 46.405 ;
      VIA 42.09 46.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 46.055 42.86 46.425 ;
      VIA 42.09 46.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 46.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 40.635 42.88 40.965 ;
      VIA 42.09 40.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 40.615 42.86 40.985 ;
      VIA 42.09 40.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 40.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 35.195 42.88 35.525 ;
      VIA 42.09 35.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 35.175 42.86 35.545 ;
      VIA 42.09 35.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 35.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 29.755 42.88 30.085 ;
      VIA 42.09 29.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 29.735 42.86 30.105 ;
      VIA 42.09 29.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 29.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 24.315 42.88 24.645 ;
      VIA 42.09 24.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 24.295 42.86 24.665 ;
      VIA 42.09 24.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 24.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 18.875 42.88 19.205 ;
      VIA 42.09 19.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 18.855 42.86 19.225 ;
      VIA 42.09 19.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 19.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 13.435 42.88 13.765 ;
      VIA 42.09 13.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 13.415 42.86 13.785 ;
      VIA 42.09 13.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 13.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 7.995 42.88 8.325 ;
      VIA 42.09 8.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 7.975 42.86 8.345 ;
      VIA 42.09 8.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 8.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  41.3 2.555 42.88 2.885 ;
      VIA 42.09 2.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  41.32 2.535 42.86 2.905 ;
      VIA 42.09 2.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 42.09 2.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 698.875 15.74 699.205 ;
      VIA 14.95 699.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 698.855 15.72 699.225 ;
      VIA 14.95 699.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 699.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 693.435 15.74 693.765 ;
      VIA 14.95 693.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 693.415 15.72 693.785 ;
      VIA 14.95 693.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 693.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 687.995 15.74 688.325 ;
      VIA 14.95 688.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 687.975 15.72 688.345 ;
      VIA 14.95 688.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 688.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 682.555 15.74 682.885 ;
      VIA 14.95 682.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 682.535 15.72 682.905 ;
      VIA 14.95 682.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 682.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 677.115 15.74 677.445 ;
      VIA 14.95 677.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 677.095 15.72 677.465 ;
      VIA 14.95 677.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 677.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 671.675 15.74 672.005 ;
      VIA 14.95 671.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 671.655 15.72 672.025 ;
      VIA 14.95 671.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 671.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 666.235 15.74 666.565 ;
      VIA 14.95 666.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 666.215 15.72 666.585 ;
      VIA 14.95 666.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 666.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 660.795 15.74 661.125 ;
      VIA 14.95 660.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 660.775 15.72 661.145 ;
      VIA 14.95 660.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 660.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 655.355 15.74 655.685 ;
      VIA 14.95 655.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 655.335 15.72 655.705 ;
      VIA 14.95 655.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 655.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 649.915 15.74 650.245 ;
      VIA 14.95 650.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 649.895 15.72 650.265 ;
      VIA 14.95 650.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 650.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 644.475 15.74 644.805 ;
      VIA 14.95 644.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 644.455 15.72 644.825 ;
      VIA 14.95 644.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 644.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 639.035 15.74 639.365 ;
      VIA 14.95 639.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 639.015 15.72 639.385 ;
      VIA 14.95 639.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 639.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 633.595 15.74 633.925 ;
      VIA 14.95 633.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 633.575 15.72 633.945 ;
      VIA 14.95 633.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 633.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 628.155 15.74 628.485 ;
      VIA 14.95 628.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 628.135 15.72 628.505 ;
      VIA 14.95 628.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 628.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 622.715 15.74 623.045 ;
      VIA 14.95 622.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 622.695 15.72 623.065 ;
      VIA 14.95 622.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 622.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 617.275 15.74 617.605 ;
      VIA 14.95 617.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 617.255 15.72 617.625 ;
      VIA 14.95 617.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 617.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 611.835 15.74 612.165 ;
      VIA 14.95 612 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 611.815 15.72 612.185 ;
      VIA 14.95 612 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 612 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 606.395 15.74 606.725 ;
      VIA 14.95 606.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 606.375 15.72 606.745 ;
      VIA 14.95 606.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 606.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 600.955 15.74 601.285 ;
      VIA 14.95 601.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 600.935 15.72 601.305 ;
      VIA 14.95 601.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 601.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 595.515 15.74 595.845 ;
      VIA 14.95 595.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 595.495 15.72 595.865 ;
      VIA 14.95 595.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 595.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 590.075 15.74 590.405 ;
      VIA 14.95 590.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 590.055 15.72 590.425 ;
      VIA 14.95 590.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 590.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 584.635 15.74 584.965 ;
      VIA 14.95 584.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 584.615 15.72 584.985 ;
      VIA 14.95 584.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 584.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 579.195 15.74 579.525 ;
      VIA 14.95 579.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 579.175 15.72 579.545 ;
      VIA 14.95 579.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 579.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 573.755 15.74 574.085 ;
      VIA 14.95 573.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 573.735 15.72 574.105 ;
      VIA 14.95 573.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 573.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 568.315 15.74 568.645 ;
      VIA 14.95 568.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 568.295 15.72 568.665 ;
      VIA 14.95 568.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 568.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 562.875 15.74 563.205 ;
      VIA 14.95 563.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 562.855 15.72 563.225 ;
      VIA 14.95 563.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 563.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 557.435 15.74 557.765 ;
      VIA 14.95 557.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 557.415 15.72 557.785 ;
      VIA 14.95 557.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 557.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 551.995 15.74 552.325 ;
      VIA 14.95 552.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 551.975 15.72 552.345 ;
      VIA 14.95 552.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 552.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 546.555 15.74 546.885 ;
      VIA 14.95 546.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 546.535 15.72 546.905 ;
      VIA 14.95 546.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 546.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 541.115 15.74 541.445 ;
      VIA 14.95 541.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 541.095 15.72 541.465 ;
      VIA 14.95 541.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 541.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 535.675 15.74 536.005 ;
      VIA 14.95 535.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 535.655 15.72 536.025 ;
      VIA 14.95 535.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 535.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 530.235 15.74 530.565 ;
      VIA 14.95 530.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 530.215 15.72 530.585 ;
      VIA 14.95 530.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 530.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 524.795 15.74 525.125 ;
      VIA 14.95 524.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 524.775 15.72 525.145 ;
      VIA 14.95 524.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 524.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 519.355 15.74 519.685 ;
      VIA 14.95 519.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 519.335 15.72 519.705 ;
      VIA 14.95 519.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 519.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 513.915 15.74 514.245 ;
      VIA 14.95 514.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 513.895 15.72 514.265 ;
      VIA 14.95 514.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 514.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 508.475 15.74 508.805 ;
      VIA 14.95 508.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 508.455 15.72 508.825 ;
      VIA 14.95 508.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 508.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 503.035 15.74 503.365 ;
      VIA 14.95 503.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 503.015 15.72 503.385 ;
      VIA 14.95 503.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 503.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 497.595 15.74 497.925 ;
      VIA 14.95 497.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 497.575 15.72 497.945 ;
      VIA 14.95 497.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 497.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 492.155 15.74 492.485 ;
      VIA 14.95 492.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 492.135 15.72 492.505 ;
      VIA 14.95 492.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 492.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 486.715 15.74 487.045 ;
      VIA 14.95 486.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 486.695 15.72 487.065 ;
      VIA 14.95 486.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 486.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 481.275 15.74 481.605 ;
      VIA 14.95 481.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 481.255 15.72 481.625 ;
      VIA 14.95 481.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 481.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 475.835 15.74 476.165 ;
      VIA 14.95 476 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 475.815 15.72 476.185 ;
      VIA 14.95 476 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 476 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 470.395 15.74 470.725 ;
      VIA 14.95 470.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 470.375 15.72 470.745 ;
      VIA 14.95 470.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 470.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 464.955 15.74 465.285 ;
      VIA 14.95 465.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 464.935 15.72 465.305 ;
      VIA 14.95 465.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 465.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 459.515 15.74 459.845 ;
      VIA 14.95 459.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 459.495 15.72 459.865 ;
      VIA 14.95 459.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 459.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 454.075 15.74 454.405 ;
      VIA 14.95 454.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 454.055 15.72 454.425 ;
      VIA 14.95 454.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 454.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 448.635 15.74 448.965 ;
      VIA 14.95 448.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 448.615 15.72 448.985 ;
      VIA 14.95 448.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 448.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 443.195 15.74 443.525 ;
      VIA 14.95 443.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 443.175 15.72 443.545 ;
      VIA 14.95 443.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 443.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 437.755 15.74 438.085 ;
      VIA 14.95 437.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 437.735 15.72 438.105 ;
      VIA 14.95 437.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 437.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 432.315 15.74 432.645 ;
      VIA 14.95 432.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 432.295 15.72 432.665 ;
      VIA 14.95 432.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 432.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 426.875 15.74 427.205 ;
      VIA 14.95 427.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 426.855 15.72 427.225 ;
      VIA 14.95 427.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 427.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 421.435 15.74 421.765 ;
      VIA 14.95 421.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 421.415 15.72 421.785 ;
      VIA 14.95 421.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 421.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 415.995 15.74 416.325 ;
      VIA 14.95 416.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 415.975 15.72 416.345 ;
      VIA 14.95 416.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 416.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 410.555 15.74 410.885 ;
      VIA 14.95 410.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 410.535 15.72 410.905 ;
      VIA 14.95 410.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 410.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 405.115 15.74 405.445 ;
      VIA 14.95 405.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 405.095 15.72 405.465 ;
      VIA 14.95 405.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 405.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 399.675 15.74 400.005 ;
      VIA 14.95 399.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 399.655 15.72 400.025 ;
      VIA 14.95 399.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 399.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 394.235 15.74 394.565 ;
      VIA 14.95 394.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 394.215 15.72 394.585 ;
      VIA 14.95 394.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 394.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 388.795 15.74 389.125 ;
      VIA 14.95 388.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 388.775 15.72 389.145 ;
      VIA 14.95 388.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 388.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 383.355 15.74 383.685 ;
      VIA 14.95 383.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 383.335 15.72 383.705 ;
      VIA 14.95 383.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 383.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 377.915 15.74 378.245 ;
      VIA 14.95 378.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 377.895 15.72 378.265 ;
      VIA 14.95 378.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 378.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 372.475 15.74 372.805 ;
      VIA 14.95 372.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 372.455 15.72 372.825 ;
      VIA 14.95 372.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 372.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 367.035 15.74 367.365 ;
      VIA 14.95 367.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 367.015 15.72 367.385 ;
      VIA 14.95 367.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 367.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 361.595 15.74 361.925 ;
      VIA 14.95 361.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 361.575 15.72 361.945 ;
      VIA 14.95 361.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 361.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 356.155 15.74 356.485 ;
      VIA 14.95 356.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 356.135 15.72 356.505 ;
      VIA 14.95 356.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 356.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 350.715 15.74 351.045 ;
      VIA 14.95 350.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 350.695 15.72 351.065 ;
      VIA 14.95 350.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 350.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 345.275 15.74 345.605 ;
      VIA 14.95 345.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 345.255 15.72 345.625 ;
      VIA 14.95 345.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 345.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 339.835 15.74 340.165 ;
      VIA 14.95 340 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 339.815 15.72 340.185 ;
      VIA 14.95 340 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 340 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 334.395 15.74 334.725 ;
      VIA 14.95 334.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 334.375 15.72 334.745 ;
      VIA 14.95 334.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 334.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 328.955 15.74 329.285 ;
      VIA 14.95 329.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 328.935 15.72 329.305 ;
      VIA 14.95 329.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 329.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 323.515 15.74 323.845 ;
      VIA 14.95 323.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 323.495 15.72 323.865 ;
      VIA 14.95 323.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 323.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 318.075 15.74 318.405 ;
      VIA 14.95 318.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 318.055 15.72 318.425 ;
      VIA 14.95 318.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 318.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 312.635 15.74 312.965 ;
      VIA 14.95 312.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 312.615 15.72 312.985 ;
      VIA 14.95 312.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 312.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 307.195 15.74 307.525 ;
      VIA 14.95 307.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 307.175 15.72 307.545 ;
      VIA 14.95 307.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 307.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 301.755 15.74 302.085 ;
      VIA 14.95 301.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 301.735 15.72 302.105 ;
      VIA 14.95 301.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 301.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 296.315 15.74 296.645 ;
      VIA 14.95 296.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 296.295 15.72 296.665 ;
      VIA 14.95 296.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 296.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 290.875 15.74 291.205 ;
      VIA 14.95 291.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 290.855 15.72 291.225 ;
      VIA 14.95 291.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 291.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 285.435 15.74 285.765 ;
      VIA 14.95 285.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 285.415 15.72 285.785 ;
      VIA 14.95 285.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 285.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 279.995 15.74 280.325 ;
      VIA 14.95 280.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 279.975 15.72 280.345 ;
      VIA 14.95 280.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 280.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 274.555 15.74 274.885 ;
      VIA 14.95 274.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 274.535 15.72 274.905 ;
      VIA 14.95 274.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 274.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 269.115 15.74 269.445 ;
      VIA 14.95 269.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 269.095 15.72 269.465 ;
      VIA 14.95 269.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 269.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 263.675 15.74 264.005 ;
      VIA 14.95 263.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 263.655 15.72 264.025 ;
      VIA 14.95 263.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 263.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 258.235 15.74 258.565 ;
      VIA 14.95 258.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 258.215 15.72 258.585 ;
      VIA 14.95 258.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 258.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 252.795 15.74 253.125 ;
      VIA 14.95 252.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 252.775 15.72 253.145 ;
      VIA 14.95 252.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 252.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 247.355 15.74 247.685 ;
      VIA 14.95 247.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 247.335 15.72 247.705 ;
      VIA 14.95 247.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 247.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 241.915 15.74 242.245 ;
      VIA 14.95 242.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 241.895 15.72 242.265 ;
      VIA 14.95 242.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 242.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 236.475 15.74 236.805 ;
      VIA 14.95 236.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 236.455 15.72 236.825 ;
      VIA 14.95 236.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 236.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 231.035 15.74 231.365 ;
      VIA 14.95 231.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 231.015 15.72 231.385 ;
      VIA 14.95 231.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 231.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 225.595 15.74 225.925 ;
      VIA 14.95 225.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 225.575 15.72 225.945 ;
      VIA 14.95 225.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 225.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 220.155 15.74 220.485 ;
      VIA 14.95 220.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 220.135 15.72 220.505 ;
      VIA 14.95 220.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 220.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 214.715 15.74 215.045 ;
      VIA 14.95 214.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 214.695 15.72 215.065 ;
      VIA 14.95 214.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 214.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 209.275 15.74 209.605 ;
      VIA 14.95 209.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 209.255 15.72 209.625 ;
      VIA 14.95 209.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 209.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 203.835 15.74 204.165 ;
      VIA 14.95 204 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 203.815 15.72 204.185 ;
      VIA 14.95 204 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 204 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 198.395 15.74 198.725 ;
      VIA 14.95 198.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 198.375 15.72 198.745 ;
      VIA 14.95 198.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 198.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 192.955 15.74 193.285 ;
      VIA 14.95 193.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 192.935 15.72 193.305 ;
      VIA 14.95 193.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 193.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 187.515 15.74 187.845 ;
      VIA 14.95 187.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 187.495 15.72 187.865 ;
      VIA 14.95 187.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 187.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 182.075 15.74 182.405 ;
      VIA 14.95 182.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 182.055 15.72 182.425 ;
      VIA 14.95 182.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 182.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 176.635 15.74 176.965 ;
      VIA 14.95 176.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 176.615 15.72 176.985 ;
      VIA 14.95 176.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 176.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 171.195 15.74 171.525 ;
      VIA 14.95 171.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 171.175 15.72 171.545 ;
      VIA 14.95 171.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 171.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 165.755 15.74 166.085 ;
      VIA 14.95 165.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 165.735 15.72 166.105 ;
      VIA 14.95 165.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 165.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 160.315 15.74 160.645 ;
      VIA 14.95 160.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 160.295 15.72 160.665 ;
      VIA 14.95 160.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 160.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 154.875 15.74 155.205 ;
      VIA 14.95 155.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 154.855 15.72 155.225 ;
      VIA 14.95 155.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 155.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 149.435 15.74 149.765 ;
      VIA 14.95 149.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 149.415 15.72 149.785 ;
      VIA 14.95 149.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 149.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 143.995 15.74 144.325 ;
      VIA 14.95 144.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 143.975 15.72 144.345 ;
      VIA 14.95 144.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 144.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 138.555 15.74 138.885 ;
      VIA 14.95 138.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 138.535 15.72 138.905 ;
      VIA 14.95 138.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 138.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 133.115 15.74 133.445 ;
      VIA 14.95 133.28 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 133.095 15.72 133.465 ;
      VIA 14.95 133.28 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 133.28 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 127.675 15.74 128.005 ;
      VIA 14.95 127.84 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 127.655 15.72 128.025 ;
      VIA 14.95 127.84 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 127.84 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 122.235 15.74 122.565 ;
      VIA 14.95 122.4 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 122.215 15.72 122.585 ;
      VIA 14.95 122.4 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 122.4 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 116.795 15.74 117.125 ;
      VIA 14.95 116.96 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 116.775 15.72 117.145 ;
      VIA 14.95 116.96 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 116.96 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 111.355 15.74 111.685 ;
      VIA 14.95 111.52 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 111.335 15.72 111.705 ;
      VIA 14.95 111.52 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 111.52 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 105.915 15.74 106.245 ;
      VIA 14.95 106.08 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 105.895 15.72 106.265 ;
      VIA 14.95 106.08 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 106.08 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 100.475 15.74 100.805 ;
      VIA 14.95 100.64 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 100.455 15.72 100.825 ;
      VIA 14.95 100.64 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 100.64 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 95.035 15.74 95.365 ;
      VIA 14.95 95.2 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 95.015 15.72 95.385 ;
      VIA 14.95 95.2 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 95.2 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 89.595 15.74 89.925 ;
      VIA 14.95 89.76 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 89.575 15.72 89.945 ;
      VIA 14.95 89.76 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 89.76 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 84.155 15.74 84.485 ;
      VIA 14.95 84.32 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 84.135 15.72 84.505 ;
      VIA 14.95 84.32 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 84.32 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 78.715 15.74 79.045 ;
      VIA 14.95 78.88 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 78.695 15.72 79.065 ;
      VIA 14.95 78.88 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 78.88 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 73.275 15.74 73.605 ;
      VIA 14.95 73.44 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 73.255 15.72 73.625 ;
      VIA 14.95 73.44 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 73.44 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 67.835 15.74 68.165 ;
      VIA 14.95 68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 67.815 15.72 68.185 ;
      VIA 14.95 68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 62.395 15.74 62.725 ;
      VIA 14.95 62.56 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 62.375 15.72 62.745 ;
      VIA 14.95 62.56 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 62.56 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 56.955 15.74 57.285 ;
      VIA 14.95 57.12 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 56.935 15.72 57.305 ;
      VIA 14.95 57.12 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 57.12 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 51.515 15.74 51.845 ;
      VIA 14.95 51.68 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 51.495 15.72 51.865 ;
      VIA 14.95 51.68 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 51.68 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 46.075 15.74 46.405 ;
      VIA 14.95 46.24 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 46.055 15.72 46.425 ;
      VIA 14.95 46.24 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 46.24 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 40.635 15.74 40.965 ;
      VIA 14.95 40.8 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 40.615 15.72 40.985 ;
      VIA 14.95 40.8 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 40.8 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 35.195 15.74 35.525 ;
      VIA 14.95 35.36 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 35.175 15.72 35.545 ;
      VIA 14.95 35.36 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 35.36 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 29.755 15.74 30.085 ;
      VIA 14.95 29.92 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 29.735 15.72 30.105 ;
      VIA 14.95 29.92 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 29.92 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 24.315 15.74 24.645 ;
      VIA 14.95 24.48 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 24.295 15.72 24.665 ;
      VIA 14.95 24.48 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 24.48 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 18.875 15.74 19.205 ;
      VIA 14.95 19.04 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 18.855 15.72 19.225 ;
      VIA 14.95 19.04 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 19.04 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 13.435 15.74 13.765 ;
      VIA 14.95 13.6 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 13.415 15.72 13.785 ;
      VIA 14.95 13.6 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 13.6 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 7.995 15.74 8.325 ;
      VIA 14.95 8.16 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 7.975 15.72 8.345 ;
      VIA 14.95 8.16 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 8.16 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  14.16 2.555 15.74 2.885 ;
      VIA 14.95 2.72 ibex_id_stage_via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  14.18 2.535 15.72 2.905 ;
      VIA 14.95 2.72 ibex_id_stage_via3_4_1600_480_1_4_400_400 ;
      VIA 14.95 2.72 ibex_id_stage_via2_3_1600_480_1_5_320_320 ;
    END
  END VSS
  PIN alu_operand_a_ex_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 165.43 177.52 165.73 ;
    END
  END alu_operand_a_ex_o[0]
  PIN alu_operand_a_ex_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 410.23 0.8 410.53 ;
    END
  END alu_operand_a_ex_o[10]
  PIN alu_operand_a_ex_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 436.75 0.8 437.05 ;
    END
  END alu_operand_a_ex_o[11]
  PIN alu_operand_a_ex_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 424.51 0.8 424.81 ;
    END
  END alu_operand_a_ex_o[12]
  PIN alu_operand_a_ex_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 636.67 0.8 636.97 ;
    END
  END alu_operand_a_ex_o[13]
  PIN alu_operand_a_ex_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 610.15 0.8 610.45 ;
    END
  END alu_operand_a_ex_o[14]
  PIN alu_operand_a_ex_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 373.51 0.8 373.81 ;
    END
  END alu_operand_a_ex_o[15]
  PIN alu_operand_a_ex_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 298.03 0.8 298.33 ;
    END
  END alu_operand_a_ex_o[16]
  PIN alu_operand_a_ex_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 344.95 0.8 345.25 ;
    END
  END alu_operand_a_ex_o[17]
  PIN alu_operand_a_ex_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 330.67 0.8 330.97 ;
    END
  END alu_operand_a_ex_o[18]
  PIN alu_operand_a_ex_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 328.63 0.8 328.93 ;
    END
  END alu_operand_a_ex_o[19]
  PIN alu_operand_a_ex_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 173.59 0.8 173.89 ;
    END
  END alu_operand_a_ex_o[1]
  PIN alu_operand_a_ex_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 193.99 0.8 194.29 ;
    END
  END alu_operand_a_ex_o[20]
  PIN alu_operand_a_ex_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 244.99 0.8 245.29 ;
    END
  END alu_operand_a_ex_o[21]
  PIN alu_operand_a_ex_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 8.35 0.8 8.65 ;
    END
  END alu_operand_a_ex_o[22]
  PIN alu_operand_a_ex_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 89.95 0.8 90.25 ;
    END
  END alu_operand_a_ex_o[23]
  PIN alu_operand_a_ex_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 271.51 0.8 271.81 ;
    END
  END alu_operand_a_ex_o[24]
  PIN alu_operand_a_ex_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 159.31 0.8 159.61 ;
    END
  END alu_operand_a_ex_o[25]
  PIN alu_operand_a_ex_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 142.99 0.8 143.29 ;
    END
  END alu_operand_a_ex_o[26]
  PIN alu_operand_a_ex_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 55.27 0.8 55.57 ;
    END
  END alu_operand_a_ex_o[27]
  PIN alu_operand_a_ex_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 30.79 0.8 31.09 ;
    END
  END alu_operand_a_ex_o[28]
  PIN alu_operand_a_ex_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 87.91 0.8 88.21 ;
    END
  END alu_operand_a_ex_o[29]
  PIN alu_operand_a_ex_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 169.51 0.8 169.81 ;
    END
  END alu_operand_a_ex_o[2]
  PIN alu_operand_a_ex_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 157.27 0.8 157.57 ;
    END
  END alu_operand_a_ex_o[30]
  PIN alu_operand_a_ex_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 75.67 177.52 75.97 ;
    END
  END alu_operand_a_ex_o[31]
  PIN alu_operand_a_ex_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 12.43 0.8 12.73 ;
    END
  END alu_operand_a_ex_o[3]
  PIN alu_operand_a_ex_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 183.79 0.8 184.09 ;
    END
  END alu_operand_a_ex_o[4]
  PIN alu_operand_a_ex_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 320.47 0.8 320.77 ;
    END
  END alu_operand_a_ex_o[5]
  PIN alu_operand_a_ex_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 340.87 0.8 341.17 ;
    END
  END alu_operand_a_ex_o[6]
  PIN alu_operand_a_ex_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 367.39 0.8 367.69 ;
    END
  END alu_operand_a_ex_o[7]
  PIN alu_operand_a_ex_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 397.99 0.8 398.29 ;
    END
  END alu_operand_a_ex_o[8]
  PIN alu_operand_a_ex_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 685.63 0.8 685.93 ;
    END
  END alu_operand_a_ex_o[9]
  PIN alu_operand_b_ex_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 571.39 0.8 571.69 ;
    END
  END alu_operand_b_ex_o[0]
  PIN alu_operand_b_ex_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 644.83 0.8 645.13 ;
    END
  END alu_operand_b_ex_o[10]
  PIN alu_operand_b_ex_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 563.23 0.8 563.53 ;
    END
  END alu_operand_b_ex_o[11]
  PIN alu_operand_b_ex_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 538.75 0.8 539.05 ;
    END
  END alu_operand_b_ex_o[12]
  PIN alu_operand_b_ex_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 473.47 0.8 473.77 ;
    END
  END alu_operand_b_ex_o[13]
  PIN alu_operand_b_ex_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 457.15 0.8 457.45 ;
    END
  END alu_operand_b_ex_o[14]
  PIN alu_operand_b_ex_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 471.43 0.8 471.73 ;
    END
  END alu_operand_b_ex_o[15]
  PIN alu_operand_b_ex_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 459.19 0.8 459.49 ;
    END
  END alu_operand_b_ex_o[16]
  PIN alu_operand_b_ex_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 565.27 0.8 565.57 ;
    END
  END alu_operand_b_ex_o[17]
  PIN alu_operand_b_ex_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 455.11 0.8 455.41 ;
    END
  END alu_operand_b_ex_o[18]
  PIN alu_operand_b_ex_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 475.51 0.8 475.81 ;
    END
  END alu_operand_b_ex_o[19]
  PIN alu_operand_b_ex_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 481.63 0.8 481.93 ;
    END
  END alu_operand_b_ex_o[1]
  PIN alu_operand_b_ex_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 548.95 0.8 549.25 ;
    END
  END alu_operand_b_ex_o[20]
  PIN alu_operand_b_ex_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 512.23 0.8 512.53 ;
    END
  END alu_operand_b_ex_o[21]
  PIN alu_operand_b_ex_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 522.43 0.8 522.73 ;
    END
  END alu_operand_b_ex_o[22]
  PIN alu_operand_b_ex_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 497.95 0.8 498.25 ;
    END
  END alu_operand_b_ex_o[23]
  PIN alu_operand_b_ex_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 524.47 0.8 524.77 ;
    END
  END alu_operand_b_ex_o[24]
  PIN alu_operand_b_ex_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 573.43 0.8 573.73 ;
    END
  END alu_operand_b_ex_o[25]
  PIN alu_operand_b_ex_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 577.51 0.8 577.81 ;
    END
  END alu_operand_b_ex_o[26]
  PIN alu_operand_b_ex_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 648.91 0.8 649.21 ;
    END
  END alu_operand_b_ex_o[27]
  PIN alu_operand_b_ex_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 614.23 0.8 614.53 ;
    END
  END alu_operand_b_ex_o[28]
  PIN alu_operand_b_ex_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 638.71 0.8 639.01 ;
    END
  END alu_operand_b_ex_o[29]
  PIN alu_operand_b_ex_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 434.71 0.8 435.01 ;
    END
  END alu_operand_b_ex_o[2]
  PIN alu_operand_b_ex_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 504.07 0.8 504.37 ;
    END
  END alu_operand_b_ex_o[30]
  PIN alu_operand_b_ex_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 520.39 0.8 520.69 ;
    END
  END alu_operand_b_ex_o[31]
  PIN alu_operand_b_ex_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 514.27 0.8 514.57 ;
    END
  END alu_operand_b_ex_o[3]
  PIN alu_operand_b_ex_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 506.11 0.8 506.41 ;
    END
  END alu_operand_b_ex_o[4]
  PIN alu_operand_b_ex_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 595.87 0.8 596.17 ;
    END
  END alu_operand_b_ex_o[5]
  PIN alu_operand_b_ex_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 632.59 177.52 632.89 ;
    END
  END alu_operand_b_ex_o[6]
  PIN alu_operand_b_ex_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 561.19 177.52 561.49 ;
    END
  END alu_operand_b_ex_o[7]
  PIN alu_operand_b_ex_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 581.59 0.8 581.89 ;
    END
  END alu_operand_b_ex_o[8]
  PIN alu_operand_b_ex_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 579.55 0.8 579.85 ;
    END
  END alu_operand_b_ex_o[9]
  PIN alu_operator_ex_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 147.07 177.52 147.37 ;
    END
  END alu_operator_ex_o[0]
  PIN alu_operator_ex_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 138.91 177.52 139.21 ;
    END
  END alu_operator_ex_o[1]
  PIN alu_operator_ex_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 191.95 177.52 192.25 ;
    END
  END alu_operator_ex_o[2]
  PIN alu_operator_ex_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 161.35 177.52 161.65 ;
    END
  END alu_operator_ex_o[3]
  PIN alu_operator_ex_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 106.27 177.52 106.57 ;
    END
  END alu_operator_ex_o[4]
  PIN alu_operator_ex_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 83.83 177.52 84.13 ;
    END
  END alu_operator_ex_o[5]
  PIN branch_decision_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 149.11 177.52 149.41 ;
    END
  END branch_decision_i
  PIN bt_a_operand_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 189.91 0.8 190.21 ;
    END
  END bt_a_operand_o[0]
  PIN bt_a_operand_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 175.63 0.8 175.93 ;
    END
  END bt_a_operand_o[10]
  PIN bt_a_operand_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 45.07 0.8 45.37 ;
    END
  END bt_a_operand_o[11]
  PIN bt_a_operand_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 59.35 0.8 59.65 ;
    END
  END bt_a_operand_o[12]
  PIN bt_a_operand_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 75.67 0.8 75.97 ;
    END
  END bt_a_operand_o[13]
  PIN bt_a_operand_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 232.75 0.8 233.05 ;
    END
  END bt_a_operand_o[14]
  PIN bt_a_operand_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 22.63 0.8 22.93 ;
    END
  END bt_a_operand_o[15]
  PIN bt_a_operand_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 226.63 0.8 226.93 ;
    END
  END bt_a_operand_o[16]
  PIN bt_a_operand_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 63.43 0.8 63.73 ;
    END
  END bt_a_operand_o[17]
  PIN bt_a_operand_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 77.71 0.8 78.01 ;
    END
  END bt_a_operand_o[18]
  PIN bt_a_operand_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 98.11 0.8 98.41 ;
    END
  END bt_a_operand_o[19]
  PIN bt_a_operand_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 83.83 0.8 84.13 ;
    END
  END bt_a_operand_o[1]
  PIN bt_a_operand_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 138.91 0.8 139.21 ;
    END
  END bt_a_operand_o[20]
  PIN bt_a_operand_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 51.19 0.8 51.49 ;
    END
  END bt_a_operand_o[21]
  PIN bt_a_operand_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 249.07 0.8 249.37 ;
    END
  END bt_a_operand_o[22]
  PIN bt_a_operand_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 185.83 0.8 186.13 ;
    END
  END bt_a_operand_o[23]
  PIN bt_a_operand_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 147.07 0.8 147.37 ;
    END
  END bt_a_operand_o[24]
  PIN bt_a_operand_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 218.47 0.8 218.77 ;
    END
  END bt_a_operand_o[25]
  PIN bt_a_operand_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 20.59 0.8 20.89 ;
    END
  END bt_a_operand_o[26]
  PIN bt_a_operand_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 161.35 0.8 161.65 ;
    END
  END bt_a_operand_o[27]
  PIN bt_a_operand_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 126.67 0.8 126.97 ;
    END
  END bt_a_operand_o[28]
  PIN bt_a_operand_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 67.51 0.8 67.81 ;
    END
  END bt_a_operand_o[29]
  PIN bt_a_operand_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 49.15 0.8 49.45 ;
    END
  END bt_a_operand_o[2]
  PIN bt_a_operand_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 34.87 0.8 35.17 ;
    END
  END bt_a_operand_o[30]
  PIN bt_a_operand_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 104.23 0.8 104.53 ;
    END
  END bt_a_operand_o[31]
  PIN bt_a_operand_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 47.11 0.8 47.41 ;
    END
  END bt_a_operand_o[3]
  PIN bt_a_operand_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 216.43 0.8 216.73 ;
    END
  END bt_a_operand_o[4]
  PIN bt_a_operand_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 124.63 0.8 124.93 ;
    END
  END bt_a_operand_o[5]
  PIN bt_a_operand_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 69.55 0.8 69.85 ;
    END
  END bt_a_operand_o[6]
  PIN bt_a_operand_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 85.87 0.8 86.17 ;
    END
  END bt_a_operand_o[7]
  PIN bt_a_operand_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 210.31 0.8 210.61 ;
    END
  END bt_a_operand_o[8]
  PIN bt_a_operand_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 110.35 0.8 110.65 ;
    END
  END bt_a_operand_o[9]
  PIN bt_b_operand_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 208.27 0.8 208.57 ;
    END
  END bt_b_operand_o[0]
  PIN bt_b_operand_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 120.55 0.8 120.85 ;
    END
  END bt_b_operand_o[10]
  PIN bt_b_operand_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 14.47 0.8 14.77 ;
    END
  END bt_b_operand_o[11]
  PIN bt_b_operand_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 65.47 0.8 65.77 ;
    END
  END bt_b_operand_o[12]
  PIN bt_b_operand_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 153.19 0.8 153.49 ;
    END
  END bt_b_operand_o[13]
  PIN bt_b_operand_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 118.51 0.8 118.81 ;
    END
  END bt_b_operand_o[14]
  PIN bt_b_operand_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 106.27 0.8 106.57 ;
    END
  END bt_b_operand_o[15]
  PIN bt_b_operand_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 177.67 0.8 177.97 ;
    END
  END bt_b_operand_o[16]
  PIN bt_b_operand_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 128.71 0.8 129.01 ;
    END
  END bt_b_operand_o[17]
  PIN bt_b_operand_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 114.43 0.8 114.73 ;
    END
  END bt_b_operand_o[18]
  PIN bt_b_operand_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 57.31 0.8 57.61 ;
    END
  END bt_b_operand_o[19]
  PIN bt_b_operand_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 32.83 0.8 33.13 ;
    END
  END bt_b_operand_o[1]
  PIN bt_b_operand_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 91.99 0.8 92.29 ;
    END
  END bt_b_operand_o[20]
  PIN bt_b_operand_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 136.87 0.8 137.17 ;
    END
  END bt_b_operand_o[21]
  PIN bt_b_operand_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 151.15 0.8 151.45 ;
    END
  END bt_b_operand_o[22]
  PIN bt_b_operand_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 165.43 0.8 165.73 ;
    END
  END bt_b_operand_o[23]
  PIN bt_b_operand_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 140.95 0.8 141.25 ;
    END
  END bt_b_operand_o[24]
  PIN bt_b_operand_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 187.87 0.8 188.17 ;
    END
  END bt_b_operand_o[25]
  PIN bt_b_operand_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 94.03 0.8 94.33 ;
    END
  END bt_b_operand_o[26]
  PIN bt_b_operand_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 206.23 0.8 206.53 ;
    END
  END bt_b_operand_o[27]
  PIN bt_b_operand_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 71.59 0.8 71.89 ;
    END
  END bt_b_operand_o[28]
  PIN bt_b_operand_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 214.39 0.8 214.69 ;
    END
  END bt_b_operand_o[29]
  PIN bt_b_operand_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 134.83 0.8 135.13 ;
    END
  END bt_b_operand_o[2]
  PIN bt_b_operand_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 16.51 0.8 16.81 ;
    END
  END bt_b_operand_o[30]
  PIN bt_b_operand_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 116.47 0.8 116.77 ;
    END
  END bt_b_operand_o[31]
  PIN bt_b_operand_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 191.95 0.8 192.25 ;
    END
  END bt_b_operand_o[3]
  PIN bt_b_operand_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 43.03 0.8 43.33 ;
    END
  END bt_b_operand_o[4]
  PIN bt_b_operand_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 220.51 0.8 220.81 ;
    END
  END bt_b_operand_o[5]
  PIN bt_b_operand_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 253.15 0.8 253.45 ;
    END
  END bt_b_operand_o[6]
  PIN bt_b_operand_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 200.11 0.8 200.41 ;
    END
  END bt_b_operand_o[7]
  PIN bt_b_operand_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 204.19 0.8 204.49 ;
    END
  END bt_b_operand_o[8]
  PIN bt_b_operand_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 73.63 0.8 73.93 ;
    END
  END bt_b_operand_o[9]
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 6.31 177.52 6.61 ;
    END
  END clk_i
  PIN csr_access_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 334.75 177.52 335.05 ;
    END
  END csr_access_o
  PIN csr_mstatus_mie_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 583.63 177.52 583.93 ;
    END
  END csr_mstatus_mie_i
  PIN csr_mstatus_tw_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 655.03 0.8 655.33 ;
    END
  END csr_mstatus_tw_i
  PIN csr_mtval_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 361.27 0.8 361.57 ;
    END
  END csr_mtval_o[0]
  PIN csr_mtval_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 400.03 0.8 400.33 ;
    END
  END csr_mtval_o[10]
  PIN csr_mtval_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 422.47 0.8 422.77 ;
    END
  END csr_mtval_o[11]
  PIN csr_mtval_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 406.15 0.8 406.45 ;
    END
  END csr_mtval_o[12]
  PIN csr_mtval_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 420.43 0.8 420.73 ;
    END
  END csr_mtval_o[13]
  PIN csr_mtval_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 618.31 0.8 618.61 ;
    END
  END csr_mtval_o[14]
  PIN csr_mtval_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 381.67 0.8 381.97 ;
    END
  END csr_mtval_o[15]
  PIN csr_mtval_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 310.27 0.8 310.57 ;
    END
  END csr_mtval_o[16]
  PIN csr_mtval_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 355.15 0.8 355.45 ;
    END
  END csr_mtval_o[17]
  PIN csr_mtval_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 324.55 0.8 324.85 ;
    END
  END csr_mtval_o[18]
  PIN csr_mtval_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 316.39 0.8 316.69 ;
    END
  END csr_mtval_o[19]
  PIN csr_mtval_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 222.55 0.8 222.85 ;
    END
  END csr_mtval_o[1]
  PIN csr_mtval_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 318.43 0.8 318.73 ;
    END
  END csr_mtval_o[20]
  PIN csr_mtval_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 24.67 0.8 24.97 ;
    END
  END csr_mtval_o[21]
  PIN csr_mtval_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 281.71 0.8 282.01 ;
    END
  END csr_mtval_o[22]
  PIN csr_mtval_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 238.87 0.8 239.17 ;
    END
  END csr_mtval_o[23]
  PIN csr_mtval_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 234.79 0.8 235.09 ;
    END
  END csr_mtval_o[24]
  PIN csr_mtval_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 149.11 0.8 149.41 ;
    END
  END csr_mtval_o[25]
  PIN csr_mtval_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 236.83 0.8 237.13 ;
    END
  END csr_mtval_o[26]
  PIN csr_mtval_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 261.31 0.8 261.61 ;
    END
  END csr_mtval_o[27]
  PIN csr_mtval_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 28.75 0.8 29.05 ;
    END
  END csr_mtval_o[28]
  PIN csr_mtval_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 112.39 0.8 112.69 ;
    END
  END csr_mtval_o[29]
  PIN csr_mtval_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 200.11 177.52 200.41 ;
    END
  END csr_mtval_o[2]
  PIN csr_mtval_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 145.03 0.8 145.33 ;
    END
  END csr_mtval_o[30]
  PIN csr_mtval_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 140.95 177.52 141.25 ;
    END
  END csr_mtval_o[31]
  PIN csr_mtval_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 110.35 177.52 110.65 ;
    END
  END csr_mtval_o[3]
  PIN csr_mtval_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 289.87 0.8 290.17 ;
    END
  END csr_mtval_o[4]
  PIN csr_mtval_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 322.51 0.8 322.81 ;
    END
  END csr_mtval_o[5]
  PIN csr_mtval_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 302.11 0.8 302.41 ;
    END
  END csr_mtval_o[6]
  PIN csr_mtval_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 363.31 0.8 363.61 ;
    END
  END csr_mtval_o[7]
  PIN csr_mtval_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 371.47 0.8 371.77 ;
    END
  END csr_mtval_o[8]
  PIN csr_mtval_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 555.07 0.8 555.37 ;
    END
  END csr_mtval_o[9]
  PIN csr_op_en_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 336.79 177.52 337.09 ;
    END
  END csr_op_en_o
  PIN csr_op_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 426.55 0.8 426.85 ;
    END
  END csr_op_o[0]
  PIN csr_op_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 567.31 0.8 567.61 ;
    END
  END csr_op_o[1]
  PIN csr_rdata_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 395.95 177.52 396.25 ;
    END
  END csr_rdata_i[0]
  PIN csr_rdata_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 391.87 177.52 392.17 ;
    END
  END csr_rdata_i[10]
  PIN csr_rdata_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 94.03 177.52 94.33 ;
    END
  END csr_rdata_i[11]
  PIN csr_rdata_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 183.79 177.52 184.09 ;
    END
  END csr_rdata_i[12]
  PIN csr_rdata_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 293.95 177.52 294.25 ;
    END
  END csr_rdata_i[13]
  PIN csr_rdata_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 295.99 177.52 296.29 ;
    END
  END csr_rdata_i[14]
  PIN csr_rdata_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 397.99 177.52 398.29 ;
    END
  END csr_rdata_i[15]
  PIN csr_rdata_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 312.31 177.52 312.61 ;
    END
  END csr_rdata_i[16]
  PIN csr_rdata_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 291.91 177.52 292.21 ;
    END
  END csr_rdata_i[17]
  PIN csr_rdata_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 10.39 177.52 10.69 ;
    END
  END csr_rdata_i[18]
  PIN csr_rdata_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 36.91 177.52 37.21 ;
    END
  END csr_rdata_i[19]
  PIN csr_rdata_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 330.67 177.52 330.97 ;
    END
  END csr_rdata_i[1]
  PIN csr_rdata_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 379.63 177.52 379.93 ;
    END
  END csr_rdata_i[20]
  PIN csr_rdata_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 402.07 177.52 402.37 ;
    END
  END csr_rdata_i[21]
  PIN csr_rdata_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 363.31 177.52 363.61 ;
    END
  END csr_rdata_i[22]
  PIN csr_rdata_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 383.71 177.52 384.01 ;
    END
  END csr_rdata_i[23]
  PIN csr_rdata_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 408.19 177.52 408.49 ;
    END
  END csr_rdata_i[24]
  PIN csr_rdata_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 332.71 177.52 333.01 ;
    END
  END csr_rdata_i[25]
  PIN csr_rdata_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 357.19 177.52 357.49 ;
    END
  END csr_rdata_i[26]
  PIN csr_rdata_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 49.15 177.52 49.45 ;
    END
  END csr_rdata_i[27]
  PIN csr_rdata_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 273.55 177.52 273.85 ;
    END
  END csr_rdata_i[28]
  PIN csr_rdata_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 318.43 177.52 318.73 ;
    END
  END csr_rdata_i[29]
  PIN csr_rdata_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 285.79 177.52 286.09 ;
    END
  END csr_rdata_i[2]
  PIN csr_rdata_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 314.35 177.52 314.65 ;
    END
  END csr_rdata_i[30]
  PIN csr_rdata_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 298.03 177.52 298.33 ;
    END
  END csr_rdata_i[31]
  PIN csr_rdata_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 316.39 177.52 316.69 ;
    END
  END csr_rdata_i[3]
  PIN csr_rdata_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 277.63 177.52 277.93 ;
    END
  END csr_rdata_i[4]
  PIN csr_rdata_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 204.19 177.52 204.49 ;
    END
  END csr_rdata_i[5]
  PIN csr_rdata_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 136.87 177.52 137.17 ;
    END
  END csr_rdata_i[6]
  PIN csr_rdata_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 263.35 177.52 263.65 ;
    END
  END csr_rdata_i[7]
  PIN csr_rdata_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 126.67 177.52 126.97 ;
    END
  END csr_rdata_i[8]
  PIN csr_rdata_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 134.83 177.52 135.13 ;
    END
  END csr_rdata_i[9]
  PIN csr_restore_dret_id_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 569.35 0.8 569.65 ;
    END
  END csr_restore_dret_id_o
  PIN csr_restore_mret_id_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 550.99 0.8 551.29 ;
    END
  END csr_restore_mret_id_o
  PIN csr_save_cause_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 628.51 0.8 628.81 ;
    END
  END csr_save_cause_o
  PIN csr_save_id_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 681.55 0.8 681.85 ;
    END
  END csr_save_id_o
  PIN csr_save_if_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 536.71 0.8 537.01 ;
    END
  END csr_save_if_o
  PIN csr_save_wb_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 96.07 0.8 96.37 ;
    END
  END csr_save_wb_o
  PIN ctrl_busy_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 536.71 177.52 537.01 ;
    END
  END ctrl_busy_o
  PIN data_ind_timing_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 310.27 177.52 310.57 ;
    END
  END data_ind_timing_i
  PIN debug_cause_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 475.51 177.52 475.81 ;
    END
  END debug_cause_o[0]
  PIN debug_cause_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 616.27 177.52 616.57 ;
    END
  END debug_cause_o[1]
  PIN debug_cause_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 542.83 177.52 543.13 ;
    END
  END debug_cause_o[2]
  PIN debug_csr_save_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 675.43 0.8 675.73 ;
    END
  END debug_csr_save_o
  PIN debug_ebreakm_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 679.51 0.8 679.81 ;
    END
  END debug_ebreakm_i
  PIN debug_ebreaku_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 559.15 0.8 559.45 ;
    END
  END debug_ebreaku_i
  PIN debug_mode_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 681.55 177.52 681.85 ;
    END
  END debug_mode_o
  PIN debug_req_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 512.23 177.52 512.53 ;
    END
  END debug_req_i
  PIN debug_single_step_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 506.11 177.52 506.41 ;
    END
  END debug_single_step_i
  PIN div_en_ex_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 189.91 177.52 190.21 ;
    END
  END div_en_ex_o
  PIN div_sel_ex_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 159.31 177.52 159.61 ;
    END
  END div_sel_ex_o
  PIN en_wb_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 349.03 177.52 349.33 ;
    END
  END en_wb_o
  PIN ex_valid_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 198.07 177.52 198.37 ;
    END
  END ex_valid_i
  PIN exc_cause_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 522.43 177.52 522.73 ;
    END
  END exc_cause_o[0]
  PIN exc_cause_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 626.47 0.8 626.77 ;
    END
  END exc_cause_o[1]
  PIN exc_cause_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 636.67 177.52 636.97 ;
    END
  END exc_cause_o[2]
  PIN exc_cause_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 534.67 0.8 534.97 ;
    END
  END exc_cause_o[3]
  PIN exc_cause_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 581.59 177.52 581.89 ;
    END
  END exc_cause_o[4]
  PIN exc_cause_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 575.47 0.8 575.77 ;
    END
  END exc_cause_o[5]
  PIN exc_pc_mux_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 673.39 0.8 673.69 ;
    END
  END exc_pc_mux_o[0]
  PIN exc_pc_mux_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 665.23 0.8 665.53 ;
    END
  END exc_pc_mux_o[1]
  PIN icache_inval_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 57.31 177.52 57.61 ;
    END
  END icache_inval_o
  PIN id_in_ready_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 387.79 0.8 388.09 ;
    END
  END id_in_ready_o
  PIN illegal_c_insn_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 220.51 177.52 220.81 ;
    END
  END illegal_c_insn_i
  PIN illegal_csr_insn_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 26.71 177.52 27.01 ;
    END
  END illegal_csr_insn_i
  PIN illegal_insn_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 532.63 0.8 532.93 ;
    END
  END illegal_insn_o
  PIN imd_val_d_ex_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 451.03 177.52 451.33 ;
    END
  END imd_val_d_ex_i[0]
  PIN imd_val_d_ex_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 493.87 177.52 494.17 ;
    END
  END imd_val_d_ex_i[10]
  PIN imd_val_d_ex_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 467.35 177.52 467.65 ;
    END
  END imd_val_d_ex_i[11]
  PIN imd_val_d_ex_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 393.91 177.52 394.21 ;
    END
  END imd_val_d_ex_i[12]
  PIN imd_val_d_ex_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 465.31 177.52 465.61 ;
    END
  END imd_val_d_ex_i[13]
  PIN imd_val_d_ex_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 377.59 177.52 377.89 ;
    END
  END imd_val_d_ex_i[14]
  PIN imd_val_d_ex_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 371.47 177.52 371.77 ;
    END
  END imd_val_d_ex_i[15]
  PIN imd_val_d_ex_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 381.67 177.52 381.97 ;
    END
  END imd_val_d_ex_i[16]
  PIN imd_val_d_ex_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 481.63 177.52 481.93 ;
    END
  END imd_val_d_ex_i[17]
  PIN imd_val_d_ex_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 487.75 177.52 488.05 ;
    END
  END imd_val_d_ex_i[18]
  PIN imd_val_d_ex_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 610.15 177.52 610.45 ;
    END
  END imd_val_d_ex_i[19]
  PIN imd_val_d_ex_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 622.39 177.52 622.69 ;
    END
  END imd_val_d_ex_i[1]
  PIN imd_val_d_ex_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 471.43 177.52 471.73 ;
    END
  END imd_val_d_ex_i[20]
  PIN imd_val_d_ex_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 508.15 177.52 508.45 ;
    END
  END imd_val_d_ex_i[21]
  PIN imd_val_d_ex_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 571.39 177.52 571.69 ;
    END
  END imd_val_d_ex_i[22]
  PIN imd_val_d_ex_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 585.67 177.52 585.97 ;
    END
  END imd_val_d_ex_i[23]
  PIN imd_val_d_ex_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 461.23 177.52 461.53 ;
    END
  END imd_val_d_ex_i[24]
  PIN imd_val_d_ex_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 516.31 177.52 516.61 ;
    END
  END imd_val_d_ex_i[25]
  PIN imd_val_d_ex_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 604.03 177.52 604.33 ;
    END
  END imd_val_d_ex_i[26]
  PIN imd_val_d_ex_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 699.91 177.52 700.21 ;
    END
  END imd_val_d_ex_i[27]
  PIN imd_val_d_ex_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 528.55 177.52 528.85 ;
    END
  END imd_val_d_ex_i[28]
  PIN imd_val_d_ex_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 557.11 177.52 557.41 ;
    END
  END imd_val_d_ex_i[29]
  PIN imd_val_d_ex_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 673.39 177.52 673.69 ;
    END
  END imd_val_d_ex_i[2]
  PIN imd_val_d_ex_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 473.47 177.52 473.77 ;
    END
  END imd_val_d_ex_i[30]
  PIN imd_val_d_ex_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 553.03 177.52 553.33 ;
    END
  END imd_val_d_ex_i[31]
  PIN imd_val_d_ex_i[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 679.51 177.52 679.81 ;
    END
  END imd_val_d_ex_i[32]
  PIN imd_val_d_ex_i[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 502.03 177.52 502.33 ;
    END
  END imd_val_d_ex_i[33]
  PIN imd_val_d_ex_i[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 302.11 177.52 302.41 ;
    END
  END imd_val_d_ex_i[34]
  PIN imd_val_d_ex_i[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 351.07 177.52 351.37 ;
    END
  END imd_val_d_ex_i[35]
  PIN imd_val_d_ex_i[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 344.95 177.52 345.25 ;
    END
  END imd_val_d_ex_i[36]
  PIN imd_val_d_ex_i[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 326.59 177.52 326.89 ;
    END
  END imd_val_d_ex_i[37]
  PIN imd_val_d_ex_i[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 281.71 177.52 282.01 ;
    END
  END imd_val_d_ex_i[38]
  PIN imd_val_d_ex_i[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 304.15 177.52 304.45 ;
    END
  END imd_val_d_ex_i[39]
  PIN imd_val_d_ex_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 504.07 177.52 504.37 ;
    END
  END imd_val_d_ex_i[3]
  PIN imd_val_d_ex_i[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 38.95 177.52 39.25 ;
    END
  END imd_val_d_ex_i[40]
  PIN imd_val_d_ex_i[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 328.63 177.52 328.93 ;
    END
  END imd_val_d_ex_i[41]
  PIN imd_val_d_ex_i[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 400.03 177.52 400.33 ;
    END
  END imd_val_d_ex_i[42]
  PIN imd_val_d_ex_i[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 73.63 177.52 73.93 ;
    END
  END imd_val_d_ex_i[43]
  PIN imd_val_d_ex_i[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 226.63 177.52 226.93 ;
    END
  END imd_val_d_ex_i[44]
  PIN imd_val_d_ex_i[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 249.07 177.52 249.37 ;
    END
  END imd_val_d_ex_i[45]
  PIN imd_val_d_ex_i[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 275.59 177.52 275.89 ;
    END
  END imd_val_d_ex_i[46]
  PIN imd_val_d_ex_i[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 216.43 177.52 216.73 ;
    END
  END imd_val_d_ex_i[47]
  PIN imd_val_d_ex_i[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 247.03 177.52 247.33 ;
    END
  END imd_val_d_ex_i[48]
  PIN imd_val_d_ex_i[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 238.87 177.52 239.17 ;
    END
  END imd_val_d_ex_i[49]
  PIN imd_val_d_ex_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 691.75 177.52 692.05 ;
    END
  END imd_val_d_ex_i[4]
  PIN imd_val_d_ex_i[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 187.87 177.52 188.17 ;
    END
  END imd_val_d_ex_i[50]
  PIN imd_val_d_ex_i[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 196.03 177.52 196.33 ;
    END
  END imd_val_d_ex_i[51]
  PIN imd_val_d_ex_i[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 228.67 177.52 228.97 ;
    END
  END imd_val_d_ex_i[52]
  PIN imd_val_d_ex_i[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 124.63 177.52 124.93 ;
    END
  END imd_val_d_ex_i[53]
  PIN imd_val_d_ex_i[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 153.19 177.52 153.49 ;
    END
  END imd_val_d_ex_i[54]
  PIN imd_val_d_ex_i[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 167.47 177.52 167.77 ;
    END
  END imd_val_d_ex_i[55]
  PIN imd_val_d_ex_i[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 112.39 177.52 112.69 ;
    END
  END imd_val_d_ex_i[56]
  PIN imd_val_d_ex_i[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 257.23 177.52 257.53 ;
    END
  END imd_val_d_ex_i[57]
  PIN imd_val_d_ex_i[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 251.11 177.52 251.41 ;
    END
  END imd_val_d_ex_i[58]
  PIN imd_val_d_ex_i[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 193.99 177.52 194.29 ;
    END
  END imd_val_d_ex_i[59]
  PIN imd_val_d_ex_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 469.39 177.52 469.69 ;
    END
  END imd_val_d_ex_i[5]
  PIN imd_val_d_ex_i[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 240.91 177.52 241.21 ;
    END
  END imd_val_d_ex_i[60]
  PIN imd_val_d_ex_i[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 163.39 177.52 163.69 ;
    END
  END imd_val_d_ex_i[61]
  PIN imd_val_d_ex_i[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 234.79 177.52 235.09 ;
    END
  END imd_val_d_ex_i[62]
  PIN imd_val_d_ex_i[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 242.95 177.52 243.25 ;
    END
  END imd_val_d_ex_i[63]
  PIN imd_val_d_ex_i[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 308.23 177.52 308.53 ;
    END
  END imd_val_d_ex_i[64]
  PIN imd_val_d_ex_i[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 283.75 177.52 284.05 ;
    END
  END imd_val_d_ex_i[65]
  PIN imd_val_d_ex_i[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 287.83 177.52 288.13 ;
    END
  END imd_val_d_ex_i[66]
  PIN imd_val_d_ex_i[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 267.43 177.52 267.73 ;
    END
  END imd_val_d_ex_i[67]
  PIN imd_val_d_ex_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 644.83 177.52 645.13 ;
    END
  END imd_val_d_ex_i[6]
  PIN imd_val_d_ex_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 479.59 177.52 479.89 ;
    END
  END imd_val_d_ex_i[7]
  PIN imd_val_d_ex_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 646.87 177.52 647.17 ;
    END
  END imd_val_d_ex_i[8]
  PIN imd_val_d_ex_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 524.47 177.52 524.77 ;
    END
  END imd_val_d_ex_i[9]
  PIN imd_val_q_ex_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 663.19 177.52 663.49 ;
    END
  END imd_val_q_ex_o[0]
  PIN imd_val_q_ex_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 695.83 177.52 696.13 ;
    END
  END imd_val_q_ex_o[10]
  PIN imd_val_q_ex_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 540.79 177.52 541.09 ;
    END
  END imd_val_q_ex_o[11]
  PIN imd_val_q_ex_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 404.11 177.52 404.41 ;
    END
  END imd_val_q_ex_o[12]
  PIN imd_val_q_ex_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 575.47 177.52 575.77 ;
    END
  END imd_val_q_ex_o[13]
  PIN imd_val_q_ex_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 406.15 177.52 406.45 ;
    END
  END imd_val_q_ex_o[14]
  PIN imd_val_q_ex_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 369.43 177.52 369.73 ;
    END
  END imd_val_q_ex_o[15]
  PIN imd_val_q_ex_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 375.55 177.52 375.85 ;
    END
  END imd_val_q_ex_o[16]
  PIN imd_val_q_ex_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 559.15 177.52 559.45 ;
    END
  END imd_val_q_ex_o[17]
  PIN imd_val_q_ex_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 426.55 177.52 426.85 ;
    END
  END imd_val_q_ex_o[18]
  PIN imd_val_q_ex_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 634.63 177.52 634.93 ;
    END
  END imd_val_q_ex_o[19]
  PIN imd_val_q_ex_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 606.07 177.52 606.37 ;
    END
  END imd_val_q_ex_o[1]
  PIN imd_val_q_ex_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 550.99 177.52 551.29 ;
    END
  END imd_val_q_ex_o[20]
  PIN imd_val_q_ex_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 597.91 177.52 598.21 ;
    END
  END imd_val_q_ex_o[21]
  PIN imd_val_q_ex_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 601.99 177.52 602.29 ;
    END
  END imd_val_q_ex_o[22]
  PIN imd_val_q_ex_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 689.71 177.52 690.01 ;
    END
  END imd_val_q_ex_o[23]
  PIN imd_val_q_ex_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 459.19 177.52 459.49 ;
    END
  END imd_val_q_ex_o[24]
  PIN imd_val_q_ex_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 463.27 177.52 463.57 ;
    END
  END imd_val_q_ex_o[25]
  PIN imd_val_q_ex_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 657.07 177.52 657.37 ;
    END
  END imd_val_q_ex_o[26]
  PIN imd_val_q_ex_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 544.87 177.52 545.17 ;
    END
  END imd_val_q_ex_o[27]
  PIN imd_val_q_ex_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 665.23 177.52 665.53 ;
    END
  END imd_val_q_ex_o[28]
  PIN imd_val_q_ex_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 687.67 177.52 687.97 ;
    END
  END imd_val_q_ex_o[29]
  PIN imd_val_q_ex_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 659.11 177.52 659.41 ;
    END
  END imd_val_q_ex_o[2]
  PIN imd_val_q_ex_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 628.51 177.52 628.81 ;
    END
  END imd_val_q_ex_o[30]
  PIN imd_val_q_ex_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 599.95 177.52 600.25 ;
    END
  END imd_val_q_ex_o[31]
  PIN imd_val_q_ex_o[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 618.31 177.52 618.61 ;
    END
  END imd_val_q_ex_o[32]
  PIN imd_val_q_ex_o[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 624.43 177.52 624.73 ;
    END
  END imd_val_q_ex_o[33]
  PIN imd_val_q_ex_o[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 71.59 177.52 71.89 ;
    END
  END imd_val_q_ex_o[34]
  PIN imd_val_q_ex_o[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 367.39 177.52 367.69 ;
    END
  END imd_val_q_ex_o[35]
  PIN imd_val_q_ex_o[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 361.27 177.52 361.57 ;
    END
  END imd_val_q_ex_o[36]
  PIN imd_val_q_ex_o[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 98.11 177.52 98.41 ;
    END
  END imd_val_q_ex_o[37]
  PIN imd_val_q_ex_o[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 269.47 177.52 269.77 ;
    END
  END imd_val_q_ex_o[38]
  PIN imd_val_q_ex_o[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 206.23 177.52 206.53 ;
    END
  END imd_val_q_ex_o[39]
  PIN imd_val_q_ex_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 608.11 177.52 608.41 ;
    END
  END imd_val_q_ex_o[3]
  PIN imd_val_q_ex_o[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 300.07 177.52 300.37 ;
    END
  END imd_val_q_ex_o[40]
  PIN imd_val_q_ex_o[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 8.35 177.52 8.65 ;
    END
  END imd_val_q_ex_o[41]
  PIN imd_val_q_ex_o[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 387.79 177.52 388.09 ;
    END
  END imd_val_q_ex_o[42]
  PIN imd_val_q_ex_o[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 320.47 177.52 320.77 ;
    END
  END imd_val_q_ex_o[43]
  PIN imd_val_q_ex_o[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 236.83 177.52 237.13 ;
    END
  END imd_val_q_ex_o[44]
  PIN imd_val_q_ex_o[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 255.19 177.52 255.49 ;
    END
  END imd_val_q_ex_o[45]
  PIN imd_val_q_ex_o[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 279.67 177.52 279.97 ;
    END
  END imd_val_q_ex_o[46]
  PIN imd_val_q_ex_o[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 67.51 177.52 67.81 ;
    END
  END imd_val_q_ex_o[47]
  PIN imd_val_q_ex_o[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 244.99 177.52 245.29 ;
    END
  END imd_val_q_ex_o[48]
  PIN imd_val_q_ex_o[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 69.55 177.52 69.85 ;
    END
  END imd_val_q_ex_o[49]
  PIN imd_val_q_ex_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 593.83 177.52 594.13 ;
    END
  END imd_val_q_ex_o[4]
  PIN imd_val_q_ex_o[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 79.75 177.52 80.05 ;
    END
  END imd_val_q_ex_o[50]
  PIN imd_val_q_ex_o[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 261.31 177.52 261.61 ;
    END
  END imd_val_q_ex_o[51]
  PIN imd_val_q_ex_o[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 230.71 177.52 231.01 ;
    END
  END imd_val_q_ex_o[52]
  PIN imd_val_q_ex_o[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 102.19 177.52 102.49 ;
    END
  END imd_val_q_ex_o[53]
  PIN imd_val_q_ex_o[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 202.15 177.52 202.45 ;
    END
  END imd_val_q_ex_o[54]
  PIN imd_val_q_ex_o[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 116.47 177.52 116.77 ;
    END
  END imd_val_q_ex_o[55]
  PIN imd_val_q_ex_o[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 185.83 177.52 186.13 ;
    END
  END imd_val_q_ex_o[56]
  PIN imd_val_q_ex_o[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 259.27 177.52 259.57 ;
    END
  END imd_val_q_ex_o[57]
  PIN imd_val_q_ex_o[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 253.15 177.52 253.45 ;
    END
  END imd_val_q_ex_o[58]
  PIN imd_val_q_ex_o[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 87.91 177.52 88.21 ;
    END
  END imd_val_q_ex_o[59]
  PIN imd_val_q_ex_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 650.95 177.52 651.25 ;
    END
  END imd_val_q_ex_o[5]
  PIN imd_val_q_ex_o[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 145.03 177.52 145.33 ;
    END
  END imd_val_q_ex_o[60]
  PIN imd_val_q_ex_o[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 222.55 177.52 222.85 ;
    END
  END imd_val_q_ex_o[61]
  PIN imd_val_q_ex_o[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 232.75 177.52 233.05 ;
    END
  END imd_val_q_ex_o[62]
  PIN imd_val_q_ex_o[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 130.75 177.52 131.05 ;
    END
  END imd_val_q_ex_o[63]
  PIN imd_val_q_ex_o[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 306.19 177.52 306.49 ;
    END
  END imd_val_q_ex_o[64]
  PIN imd_val_q_ex_o[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 212.35 177.52 212.65 ;
    END
  END imd_val_q_ex_o[65]
  PIN imd_val_q_ex_o[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 289.87 177.52 290.17 ;
    END
  END imd_val_q_ex_o[66]
  PIN imd_val_q_ex_o[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 265.39 177.52 265.69 ;
    END
  END imd_val_q_ex_o[67]
  PIN imd_val_q_ex_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 455.11 177.52 455.41 ;
    END
  END imd_val_q_ex_o[6]
  PIN imd_val_q_ex_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 424.51 177.52 424.81 ;
    END
  END imd_val_q_ex_o[7]
  PIN imd_val_q_ex_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 546.91 177.52 547.21 ;
    END
  END imd_val_q_ex_o[8]
  PIN imd_val_q_ex_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 483.67 177.52 483.97 ;
    END
  END imd_val_q_ex_o[9]
  PIN imd_val_we_ex_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 271.51 177.52 271.81 ;
    END
  END imd_val_we_ex_i[0]
  PIN imd_val_we_ex_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 630.55 177.52 630.85 ;
    END
  END imd_val_we_ex_i[1]
  PIN instr_bp_taken_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  9.36 0 9.5 0.485 ;
    END
  END instr_bp_taken_i
  PIN instr_fetch_err_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 353.11 177.52 353.41 ;
    END
  END instr_fetch_err_i
  PIN instr_fetch_err_plus2_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 10.39 0.8 10.69 ;
    END
  END instr_fetch_err_plus2_i
  PIN instr_first_cycle_id_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 181.75 177.52 182.05 ;
    END
  END instr_first_cycle_id_o
  PIN instr_id_done_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 342.91 177.52 343.21 ;
    END
  END instr_id_done_o
  PIN instr_is_compressed_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 693.79 0.8 694.09 ;
    END
  END instr_is_compressed_i
  PIN instr_perf_count_id_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 383.71 0.8 384.01 ;
    END
  END instr_perf_count_id_o
  PIN instr_rdata_alu_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 122.59 0.8 122.89 ;
    END
  END instr_rdata_alu_i[0]
  PIN instr_rdata_alu_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  160.24 0 160.38 0.485 ;
    END
  END instr_rdata_alu_i[10]
  PIN instr_rdata_alu_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  162.08 0 162.22 0.485 ;
    END
  END instr_rdata_alu_i[11]
  PIN instr_rdata_alu_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 151.15 177.52 151.45 ;
    END
  END instr_rdata_alu_i[12]
  PIN instr_rdata_alu_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 177.67 177.52 177.97 ;
    END
  END instr_rdata_alu_i[13]
  PIN instr_rdata_alu_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 173.59 177.52 173.89 ;
    END
  END instr_rdata_alu_i[14]
  PIN instr_rdata_alu_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  13.04 0 13.18 0.485 ;
    END
  END instr_rdata_alu_i[15]
  PIN instr_rdata_alu_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  145.52 0 145.66 0.485 ;
    END
  END instr_rdata_alu_i[16]
  PIN instr_rdata_alu_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  173.12 0 173.26 0.485 ;
    END
  END instr_rdata_alu_i[17]
  PIN instr_rdata_alu_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  158.4 0 158.54 0.485 ;
    END
  END instr_rdata_alu_i[18]
  PIN instr_rdata_alu_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  3.84 0 3.98 0.485 ;
    END
  END instr_rdata_alu_i[19]
  PIN instr_rdata_alu_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 130.75 0.8 131.05 ;
    END
  END instr_rdata_alu_i[1]
  PIN instr_rdata_alu_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  2 0 2.14 0.485 ;
    END
  END instr_rdata_alu_i[20]
  PIN instr_rdata_alu_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  71.92 0 72.06 0.485 ;
    END
  END instr_rdata_alu_i[21]
  PIN instr_rdata_alu_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  108.72 0 108.86 0.485 ;
    END
  END instr_rdata_alu_i[22]
  PIN instr_rdata_alu_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  48 0 48.14 0.485 ;
    END
  END instr_rdata_alu_i[23]
  PIN instr_rdata_alu_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  154.72 0 154.86 0.485 ;
    END
  END instr_rdata_alu_i[24]
  PIN instr_rdata_alu_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 142.99 177.52 143.29 ;
    END
  END instr_rdata_alu_i[25]
  PIN instr_rdata_alu_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 96.07 177.52 96.37 ;
    END
  END instr_rdata_alu_i[26]
  PIN instr_rdata_alu_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 155.23 0.8 155.53 ;
    END
  END instr_rdata_alu_i[27]
  PIN instr_rdata_alu_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 40.99 0.8 41.29 ;
    END
  END instr_rdata_alu_i[28]
  PIN instr_rdata_alu_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 167.47 0.8 167.77 ;
    END
  END instr_rdata_alu_i[29]
  PIN instr_rdata_alu_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 53.23 0.8 53.53 ;
    END
  END instr_rdata_alu_i[2]
  PIN instr_rdata_alu_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 114.43 177.52 114.73 ;
    END
  END instr_rdata_alu_i[30]
  PIN instr_rdata_alu_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 81.79 0.8 82.09 ;
    END
  END instr_rdata_alu_i[31]
  PIN instr_rdata_alu_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 132.79 0.8 133.09 ;
    END
  END instr_rdata_alu_i[3]
  PIN instr_rdata_alu_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 104.23 177.52 104.53 ;
    END
  END instr_rdata_alu_i[4]
  PIN instr_rdata_alu_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 118.51 177.52 118.81 ;
    END
  END instr_rdata_alu_i[5]
  PIN instr_rdata_alu_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 163.39 0.8 163.69 ;
    END
  END instr_rdata_alu_i[6]
  PIN instr_rdata_alu_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  152.88 0 153.02 0.485 ;
    END
  END instr_rdata_alu_i[7]
  PIN instr_rdata_alu_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  143.68 0 143.82 0.485 ;
    END
  END instr_rdata_alu_i[8]
  PIN instr_rdata_alu_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  5.68 0 5.82 0.485 ;
    END
  END instr_rdata_alu_i[9]
  PIN instr_rdata_c_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 353.11 0.8 353.41 ;
    END
  END instr_rdata_c_i[0]
  PIN instr_rdata_c_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 530.59 0.8 530.89 ;
    END
  END instr_rdata_c_i[10]
  PIN instr_rdata_c_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 430.63 0.8 430.93 ;
    END
  END instr_rdata_c_i[11]
  PIN instr_rdata_c_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 418.39 0.8 418.69 ;
    END
  END instr_rdata_c_i[12]
  PIN instr_rdata_c_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 597.91 0.8 598.21 ;
    END
  END instr_rdata_c_i[13]
  PIN instr_rdata_c_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 393.91 0.8 394.21 ;
    END
  END instr_rdata_c_i[14]
  PIN instr_rdata_c_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 379.63 0.8 379.93 ;
    END
  END instr_rdata_c_i[15]
  PIN instr_rdata_c_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 28.75 177.52 29.05 ;
    END
  END instr_rdata_c_i[1]
  PIN instr_rdata_c_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 24.67 177.52 24.97 ;
    END
  END instr_rdata_c_i[2]
  PIN instr_rdata_c_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 81.79 177.52 82.09 ;
    END
  END instr_rdata_c_i[3]
  PIN instr_rdata_c_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 14.47 177.52 14.77 ;
    END
  END instr_rdata_c_i[4]
  PIN instr_rdata_c_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 40.99 177.52 41.29 ;
    END
  END instr_rdata_c_i[5]
  PIN instr_rdata_c_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 332.71 0.8 333.01 ;
    END
  END instr_rdata_c_i[6]
  PIN instr_rdata_c_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 404.11 0.8 404.41 ;
    END
  END instr_rdata_c_i[7]
  PIN instr_rdata_c_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 412.27 0.8 412.57 ;
    END
  END instr_rdata_c_i[8]
  PIN instr_rdata_c_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 385.75 0.8 386.05 ;
    END
  END instr_rdata_c_i[9]
  PIN instr_rdata_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 4.27 177.52 4.57 ;
    END
  END instr_rdata_i[0]
  PIN instr_rdata_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 642.79 0.8 643.09 ;
    END
  END instr_rdata_i[10]
  PIN instr_rdata_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 650.95 0.8 651.25 ;
    END
  END instr_rdata_i[11]
  PIN instr_rdata_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 340.87 177.52 341.17 ;
    END
  END instr_rdata_i[12]
  PIN instr_rdata_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 338.83 0.8 339.13 ;
    END
  END instr_rdata_i[13]
  PIN instr_rdata_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 300.07 0.8 300.37 ;
    END
  END instr_rdata_i[14]
  PIN instr_rdata_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 557.11 0.8 557.41 ;
    END
  END instr_rdata_i[15]
  PIN instr_rdata_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 295.99 0.8 296.29 ;
    END
  END instr_rdata_i[16]
  PIN instr_rdata_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 293.95 0.8 294.25 ;
    END
  END instr_rdata_i[17]
  PIN instr_rdata_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 306.19 0.8 306.49 ;
    END
  END instr_rdata_i[18]
  PIN instr_rdata_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 663.19 0.8 663.49 ;
    END
  END instr_rdata_i[19]
  PIN instr_rdata_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 55.27 177.52 55.57 ;
    END
  END instr_rdata_i[1]
  PIN instr_rdata_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 683.59 0.8 683.89 ;
    END
  END instr_rdata_i[20]
  PIN instr_rdata_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 691.75 0.8 692.05 ;
    END
  END instr_rdata_i[21]
  PIN instr_rdata_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 661.15 0.8 661.45 ;
    END
  END instr_rdata_i[22]
  PIN instr_rdata_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 697.87 0.8 698.17 ;
    END
  END instr_rdata_i[23]
  PIN instr_rdata_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 695.83 0.8 696.13 ;
    END
  END instr_rdata_i[24]
  PIN instr_rdata_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 606.07 0.8 606.37 ;
    END
  END instr_rdata_i[25]
  PIN instr_rdata_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 624.43 0.8 624.73 ;
    END
  END instr_rdata_i[26]
  PIN instr_rdata_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 689.71 0.8 690.01 ;
    END
  END instr_rdata_i[27]
  PIN instr_rdata_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 699.91 0.8 700.21 ;
    END
  END instr_rdata_i[28]
  PIN instr_rdata_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 687.67 0.8 687.97 ;
    END
  END instr_rdata_i[29]
  PIN instr_rdata_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 61.39 177.52 61.69 ;
    END
  END instr_rdata_i[2]
  PIN instr_rdata_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 604.03 0.8 604.33 ;
    END
  END instr_rdata_i[30]
  PIN instr_rdata_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 585.67 0.8 585.97 ;
    END
  END instr_rdata_i[31]
  PIN instr_rdata_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 51.19 177.52 51.49 ;
    END
  END instr_rdata_i[3]
  PIN instr_rdata_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 85.87 177.52 86.17 ;
    END
  END instr_rdata_i[4]
  PIN instr_rdata_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 22.63 177.52 22.93 ;
    END
  END instr_rdata_i[5]
  PIN instr_rdata_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 157.27 177.52 157.57 ;
    END
  END instr_rdata_i[6]
  PIN instr_rdata_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 671.35 0.8 671.65 ;
    END
  END instr_rdata_i[7]
  PIN instr_rdata_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 542.83 0.8 543.13 ;
    END
  END instr_rdata_i[8]
  PIN instr_rdata_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 553.03 0.8 553.33 ;
    END
  END instr_rdata_i[9]
  PIN instr_req_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 675.43 177.52 675.73 ;
    END
  END instr_req_o
  PIN instr_type_wb_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 26.71 0.8 27.01 ;
    END
  END instr_type_wb_o[0]
  PIN instr_type_wb_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 428.59 0.8 428.89 ;
    END
  END instr_type_wb_o[1]
  PIN instr_valid_clear_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 634.63 0.8 634.93 ;
    END
  END instr_valid_clear_o
  PIN instr_valid_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 65.47 177.52 65.77 ;
    END
  END instr_valid_i
  PIN irq_nm_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 685.63 177.52 685.93 ;
    END
  END irq_nm_i
  PIN irq_pending_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 661.15 177.52 661.45 ;
    END
  END irq_pending_i
  PIN irqs_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 532.63 177.52 532.93 ;
    END
  END irqs_i[0]
  PIN irqs_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 548.95 177.52 549.25 ;
    END
  END irqs_i[10]
  PIN irqs_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 677.47 177.52 677.77 ;
    END
  END irqs_i[11]
  PIN irqs_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 589.75 177.52 590.05 ;
    END
  END irqs_i[12]
  PIN irqs_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 693.79 177.52 694.09 ;
    END
  END irqs_i[13]
  PIN irqs_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 530.59 177.52 530.89 ;
    END
  END irqs_i[14]
  PIN irqs_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 579.55 177.52 579.85 ;
    END
  END irqs_i[15]
  PIN irqs_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  94 0 94.14 0.485 ;
    END
  END irqs_i[16]
  PIN irqs_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 563.23 177.52 563.53 ;
    END
  END irqs_i[17]
  PIN irqs_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 671.35 177.52 671.65 ;
    END
  END irqs_i[1]
  PIN irqs_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 591.79 177.52 592.09 ;
    END
  END irqs_i[2]
  PIN irqs_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 569.35 177.52 569.65 ;
    END
  END irqs_i[3]
  PIN irqs_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 577.51 177.52 577.81 ;
    END
  END irqs_i[4]
  PIN irqs_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 626.47 177.52 626.77 ;
    END
  END irqs_i[5]
  PIN irqs_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 567.31 177.52 567.61 ;
    END
  END irqs_i[6]
  PIN irqs_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 655.03 177.52 655.33 ;
    END
  END irqs_i[7]
  PIN irqs_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 669.31 177.52 669.61 ;
    END
  END irqs_i[8]
  PIN irqs_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 565.27 177.52 565.57 ;
    END
  END irqs_i[9]
  PIN lsu_addr_incr_req_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 53.23 177.52 53.53 ;
    END
  END lsu_addr_incr_req_i
  PIN lsu_addr_last_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 359.23 0.8 359.53 ;
    END
  END lsu_addr_last_i[0]
  PIN lsu_addr_last_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 612.19 0.8 612.49 ;
    END
  END lsu_addr_last_i[10]
  PIN lsu_addr_last_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 432.67 0.8 432.97 ;
    END
  END lsu_addr_last_i[11]
  PIN lsu_addr_last_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 414.31 0.8 414.61 ;
    END
  END lsu_addr_last_i[12]
  PIN lsu_addr_last_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 446.95 0.8 447.25 ;
    END
  END lsu_addr_last_i[13]
  PIN lsu_addr_last_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 632.59 0.8 632.89 ;
    END
  END lsu_addr_last_i[14]
  PIN lsu_addr_last_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 377.59 0.8 377.89 ;
    END
  END lsu_addr_last_i[15]
  PIN lsu_addr_last_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 349.03 0.8 349.33 ;
    END
  END lsu_addr_last_i[16]
  PIN lsu_addr_last_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 357.19 0.8 357.49 ;
    END
  END lsu_addr_last_i[17]
  PIN lsu_addr_last_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 336.79 0.8 337.09 ;
    END
  END lsu_addr_last_i[18]
  PIN lsu_addr_last_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 334.75 0.8 335.05 ;
    END
  END lsu_addr_last_i[19]
  PIN lsu_addr_last_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 100.15 0.8 100.45 ;
    END
  END lsu_addr_last_i[1]
  PIN lsu_addr_last_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 275.59 0.8 275.89 ;
    END
  END lsu_addr_last_i[20]
  PIN lsu_addr_last_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 255.19 0.8 255.49 ;
    END
  END lsu_addr_last_i[21]
  PIN lsu_addr_last_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 269.47 0.8 269.77 ;
    END
  END lsu_addr_last_i[22]
  PIN lsu_addr_last_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 267.43 0.8 267.73 ;
    END
  END lsu_addr_last_i[23]
  PIN lsu_addr_last_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 247.03 0.8 247.33 ;
    END
  END lsu_addr_last_i[24]
  PIN lsu_addr_last_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 230.71 0.8 231.01 ;
    END
  END lsu_addr_last_i[25]
  PIN lsu_addr_last_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 224.59 0.8 224.89 ;
    END
  END lsu_addr_last_i[26]
  PIN lsu_addr_last_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 202.15 0.8 202.45 ;
    END
  END lsu_addr_last_i[27]
  PIN lsu_addr_last_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 181.75 0.8 182.05 ;
    END
  END lsu_addr_last_i[28]
  PIN lsu_addr_last_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 4.27 0.8 4.57 ;
    END
  END lsu_addr_last_i[29]
  PIN lsu_addr_last_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 32.83 177.52 33.13 ;
    END
  END lsu_addr_last_i[2]
  PIN lsu_addr_last_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 89.95 177.52 90.25 ;
    END
  END lsu_addr_last_i[30]
  PIN lsu_addr_last_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 30.79 177.52 31.09 ;
    END
  END lsu_addr_last_i[31]
  PIN lsu_addr_last_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 77.71 177.52 78.01 ;
    END
  END lsu_addr_last_i[3]
  PIN lsu_addr_last_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 314.35 0.8 314.65 ;
    END
  END lsu_addr_last_i[4]
  PIN lsu_addr_last_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 12.43 177.52 12.73 ;
    END
  END lsu_addr_last_i[5]
  PIN lsu_addr_last_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 342.91 0.8 343.21 ;
    END
  END lsu_addr_last_i[6]
  PIN lsu_addr_last_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 369.43 0.8 369.73 ;
    END
  END lsu_addr_last_i[7]
  PIN lsu_addr_last_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 659.11 0.8 659.41 ;
    END
  END lsu_addr_last_i[8]
  PIN lsu_addr_last_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 391.87 0.8 392.17 ;
    END
  END lsu_addr_last_i[9]
  PIN lsu_load_err_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 677.47 0.8 677.77 ;
    END
  END lsu_load_err_i
  PIN lsu_req_done_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  75.6 0 75.74 0.485 ;
    END
  END lsu_req_done_i
  PIN lsu_req_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 169.51 177.52 169.81 ;
    END
  END lsu_req_o
  PIN lsu_resp_valid_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 59.35 177.52 59.65 ;
    END
  END lsu_resp_valid_i
  PIN lsu_sign_ext_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 359.23 177.52 359.53 ;
    END
  END lsu_sign_ext_o
  PIN lsu_store_err_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 616.27 0.8 616.57 ;
    END
  END lsu_store_err_i
  PIN lsu_type_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 351.07 0.8 351.37 ;
    END
  END lsu_type_o[0]
  PIN lsu_type_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 355.15 177.52 355.45 ;
    END
  END lsu_type_o[1]
  PIN lsu_wdata_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 589.75 0.8 590.05 ;
    END
  END lsu_wdata_o[0]
  PIN lsu_wdata_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 640.75 0.8 641.05 ;
    END
  END lsu_wdata_o[10]
  PIN lsu_wdata_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 451.03 0.8 451.33 ;
    END
  END lsu_wdata_o[11]
  PIN lsu_wdata_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 467.35 0.8 467.65 ;
    END
  END lsu_wdata_o[12]
  PIN lsu_wdata_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 491.83 0.8 492.13 ;
    END
  END lsu_wdata_o[13]
  PIN lsu_wdata_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 463.27 0.8 463.57 ;
    END
  END lsu_wdata_o[14]
  PIN lsu_wdata_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 479.59 0.8 479.89 ;
    END
  END lsu_wdata_o[15]
  PIN lsu_wdata_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 593.83 0.8 594.13 ;
    END
  END lsu_wdata_o[16]
  PIN lsu_wdata_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 493.87 0.8 494.17 ;
    END
  END lsu_wdata_o[17]
  PIN lsu_wdata_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 453.07 0.8 453.37 ;
    END
  END lsu_wdata_o[18]
  PIN lsu_wdata_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 483.67 0.8 483.97 ;
    END
  END lsu_wdata_o[19]
  PIN lsu_wdata_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 487.75 0.8 488.05 ;
    END
  END lsu_wdata_o[1]
  PIN lsu_wdata_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 587.71 0.8 588.01 ;
    END
  END lsu_wdata_o[20]
  PIN lsu_wdata_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 561.19 0.8 561.49 ;
    END
  END lsu_wdata_o[21]
  PIN lsu_wdata_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 599.95 0.8 600.25 ;
    END
  END lsu_wdata_o[22]
  PIN lsu_wdata_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 502.03 0.8 502.33 ;
    END
  END lsu_wdata_o[23]
  PIN lsu_wdata_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 622.39 0.8 622.69 ;
    END
  END lsu_wdata_o[24]
  PIN lsu_wdata_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 642.79 177.52 643.09 ;
    END
  END lsu_wdata_o[25]
  PIN lsu_wdata_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 612.19 177.52 612.49 ;
    END
  END lsu_wdata_o[26]
  PIN lsu_wdata_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 546.91 0.8 547.21 ;
    END
  END lsu_wdata_o[27]
  PIN lsu_wdata_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 526.51 0.8 526.81 ;
    END
  END lsu_wdata_o[28]
  PIN lsu_wdata_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 508.15 0.8 508.45 ;
    END
  END lsu_wdata_o[29]
  PIN lsu_wdata_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 442.87 0.8 443.17 ;
    END
  END lsu_wdata_o[2]
  PIN lsu_wdata_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 620.35 0.8 620.65 ;
    END
  END lsu_wdata_o[30]
  PIN lsu_wdata_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 657.07 0.8 657.37 ;
    END
  END lsu_wdata_o[31]
  PIN lsu_wdata_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 518.35 0.8 518.65 ;
    END
  END lsu_wdata_o[3]
  PIN lsu_wdata_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 495.91 0.8 496.21 ;
    END
  END lsu_wdata_o[4]
  PIN lsu_wdata_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 595.87 177.52 596.17 ;
    END
  END lsu_wdata_o[5]
  PIN lsu_wdata_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 555.07 177.52 555.37 ;
    END
  END lsu_wdata_o[6]
  PIN lsu_wdata_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 587.71 177.52 588.01 ;
    END
  END lsu_wdata_o[7]
  PIN lsu_wdata_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 652.99 0.8 653.29 ;
    END
  END lsu_wdata_o[8]
  PIN lsu_wdata_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 544.87 0.8 545.17 ;
    END
  END lsu_wdata_o[9]
  PIN lsu_we_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 47.11 177.52 47.41 ;
    END
  END lsu_we_o
  PIN mult_en_ex_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 132.79 177.52 133.09 ;
    END
  END mult_en_ex_o
  PIN mult_sel_ex_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 155.23 177.52 155.53 ;
    END
  END mult_sel_ex_o
  PIN multdiv_operand_a_ex_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 100.15 177.52 100.45 ;
    END
  END multdiv_operand_a_ex_o[0]
  PIN multdiv_operand_a_ex_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 408.19 0.8 408.49 ;
    END
  END multdiv_operand_a_ex_o[10]
  PIN multdiv_operand_a_ex_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 444.91 0.8 445.21 ;
    END
  END multdiv_operand_a_ex_o[11]
  PIN multdiv_operand_a_ex_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 416.35 0.8 416.65 ;
    END
  END multdiv_operand_a_ex_o[12]
  PIN multdiv_operand_a_ex_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 438.79 0.8 439.09 ;
    END
  END multdiv_operand_a_ex_o[13]
  PIN multdiv_operand_a_ex_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 395.95 0.8 396.25 ;
    END
  END multdiv_operand_a_ex_o[14]
  PIN multdiv_operand_a_ex_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 375.55 0.8 375.85 ;
    END
  END multdiv_operand_a_ex_o[15]
  PIN multdiv_operand_a_ex_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 304.15 0.8 304.45 ;
    END
  END multdiv_operand_a_ex_o[16]
  PIN multdiv_operand_a_ex_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 312.31 0.8 312.61 ;
    END
  END multdiv_operand_a_ex_o[17]
  PIN multdiv_operand_a_ex_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 308.23 0.8 308.53 ;
    END
  END multdiv_operand_a_ex_o[18]
  PIN multdiv_operand_a_ex_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 326.59 0.8 326.89 ;
    END
  END multdiv_operand_a_ex_o[19]
  PIN multdiv_operand_a_ex_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 179.71 0.8 180.01 ;
    END
  END multdiv_operand_a_ex_o[1]
  PIN multdiv_operand_a_ex_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 277.63 0.8 277.93 ;
    END
  END multdiv_operand_a_ex_o[20]
  PIN multdiv_operand_a_ex_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 265.39 0.8 265.69 ;
    END
  END multdiv_operand_a_ex_o[21]
  PIN multdiv_operand_a_ex_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 263.35 0.8 263.65 ;
    END
  END multdiv_operand_a_ex_o[22]
  PIN multdiv_operand_a_ex_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 251.11 0.8 251.41 ;
    END
  END multdiv_operand_a_ex_o[23]
  PIN multdiv_operand_a_ex_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 36.91 0.8 37.21 ;
    END
  END multdiv_operand_a_ex_o[24]
  PIN multdiv_operand_a_ex_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 228.67 0.8 228.97 ;
    END
  END multdiv_operand_a_ex_o[25]
  PIN multdiv_operand_a_ex_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 102.19 0.8 102.49 ;
    END
  END multdiv_operand_a_ex_o[26]
  PIN multdiv_operand_a_ex_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 212.35 0.8 212.65 ;
    END
  END multdiv_operand_a_ex_o[27]
  PIN multdiv_operand_a_ex_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 61.39 0.8 61.69 ;
    END
  END multdiv_operand_a_ex_o[28]
  PIN multdiv_operand_a_ex_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 38.95 0.8 39.25 ;
    END
  END multdiv_operand_a_ex_o[29]
  PIN multdiv_operand_a_ex_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 108.31 0.8 108.61 ;
    END
  END multdiv_operand_a_ex_o[2]
  PIN multdiv_operand_a_ex_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 108.31 177.52 108.61 ;
    END
  END multdiv_operand_a_ex_o[30]
  PIN multdiv_operand_a_ex_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 218.47 177.52 218.77 ;
    END
  END multdiv_operand_a_ex_o[31]
  PIN multdiv_operand_a_ex_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 196.03 0.8 196.33 ;
    END
  END multdiv_operand_a_ex_o[3]
  PIN multdiv_operand_a_ex_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 171.55 0.8 171.85 ;
    END
  END multdiv_operand_a_ex_o[4]
  PIN multdiv_operand_a_ex_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 18.55 177.52 18.85 ;
    END
  END multdiv_operand_a_ex_o[5]
  PIN multdiv_operand_a_ex_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 346.99 0.8 347.29 ;
    END
  END multdiv_operand_a_ex_o[6]
  PIN multdiv_operand_a_ex_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 365.35 0.8 365.65 ;
    END
  END multdiv_operand_a_ex_o[7]
  PIN multdiv_operand_a_ex_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 402.07 0.8 402.37 ;
    END
  END multdiv_operand_a_ex_o[8]
  PIN multdiv_operand_a_ex_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 389.83 0.8 390.13 ;
    END
  END multdiv_operand_a_ex_o[9]
  PIN multdiv_operand_b_ex_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 669.31 0.8 669.61 ;
    END
  END multdiv_operand_b_ex_o[0]
  PIN multdiv_operand_b_ex_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 583.63 0.8 583.93 ;
    END
  END multdiv_operand_b_ex_o[10]
  PIN multdiv_operand_b_ex_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 448.99 0.8 449.29 ;
    END
  END multdiv_operand_b_ex_o[11]
  PIN multdiv_operand_b_ex_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 469.39 0.8 469.69 ;
    END
  END multdiv_operand_b_ex_o[12]
  PIN multdiv_operand_b_ex_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 489.79 0.8 490.09 ;
    END
  END multdiv_operand_b_ex_o[13]
  PIN multdiv_operand_b_ex_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 461.23 0.8 461.53 ;
    END
  END multdiv_operand_b_ex_o[14]
  PIN multdiv_operand_b_ex_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 477.55 0.8 477.85 ;
    END
  END multdiv_operand_b_ex_o[15]
  PIN multdiv_operand_b_ex_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 465.31 0.8 465.61 ;
    END
  END multdiv_operand_b_ex_o[16]
  PIN multdiv_operand_b_ex_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 630.55 0.8 630.85 ;
    END
  END multdiv_operand_b_ex_o[17]
  PIN multdiv_operand_b_ex_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 591.79 0.8 592.09 ;
    END
  END multdiv_operand_b_ex_o[18]
  PIN multdiv_operand_b_ex_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 485.71 0.8 486.01 ;
    END
  END multdiv_operand_b_ex_o[19]
  PIN multdiv_operand_b_ex_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 646.87 0.8 647.17 ;
    END
  END multdiv_operand_b_ex_o[1]
  PIN multdiv_operand_b_ex_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 667.27 0.8 667.57 ;
    END
  END multdiv_operand_b_ex_o[20]
  PIN multdiv_operand_b_ex_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 516.31 0.8 516.61 ;
    END
  END multdiv_operand_b_ex_o[21]
  PIN multdiv_operand_b_ex_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 540.79 0.8 541.09 ;
    END
  END multdiv_operand_b_ex_o[22]
  PIN multdiv_operand_b_ex_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 499.99 0.8 500.29 ;
    END
  END multdiv_operand_b_ex_o[23]
  PIN multdiv_operand_b_ex_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 608.11 0.8 608.41 ;
    END
  END multdiv_operand_b_ex_o[24]
  PIN multdiv_operand_b_ex_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 652.99 177.52 653.29 ;
    END
  END multdiv_operand_b_ex_o[25]
  PIN multdiv_operand_b_ex_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 640.75 177.52 641.05 ;
    END
  END multdiv_operand_b_ex_o[26]
  PIN multdiv_operand_b_ex_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 601.99 0.8 602.29 ;
    END
  END multdiv_operand_b_ex_o[27]
  PIN multdiv_operand_b_ex_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 528.55 0.8 528.85 ;
    END
  END multdiv_operand_b_ex_o[28]
  PIN multdiv_operand_b_ex_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 510.19 0.8 510.49 ;
    END
  END multdiv_operand_b_ex_o[29]
  PIN multdiv_operand_b_ex_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 440.83 0.8 441.13 ;
    END
  END multdiv_operand_b_ex_o[2]
  PIN multdiv_operand_b_ex_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 499.99 177.52 500.29 ;
    END
  END multdiv_operand_b_ex_o[30]
  PIN multdiv_operand_b_ex_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 683.59 177.52 683.89 ;
    END
  END multdiv_operand_b_ex_o[31]
  PIN multdiv_operand_b_ex_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 534.67 177.52 534.97 ;
    END
  END multdiv_operand_b_ex_o[3]
  PIN multdiv_operand_b_ex_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 667.27 177.52 667.57 ;
    END
  END multdiv_operand_b_ex_o[4]
  PIN multdiv_operand_b_ex_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 638.71 177.52 639.01 ;
    END
  END multdiv_operand_b_ex_o[5]
  PIN multdiv_operand_b_ex_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 620.35 177.52 620.65 ;
    END
  END multdiv_operand_b_ex_o[6]
  PIN multdiv_operand_b_ex_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 573.43 177.52 573.73 ;
    END
  END multdiv_operand_b_ex_o[7]
  PIN multdiv_operand_b_ex_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 520.39 177.52 520.69 ;
    END
  END multdiv_operand_b_ex_o[8]
  PIN multdiv_operand_b_ex_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 510.19 177.52 510.49 ;
    END
  END multdiv_operand_b_ex_o[9]
  PIN multdiv_operator_ex_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 416.35 177.52 416.65 ;
    END
  END multdiv_operator_ex_o[0]
  PIN multdiv_operator_ex_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 436.75 177.52 437.05 ;
    END
  END multdiv_operator_ex_o[1]
  PIN multdiv_ready_id_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 122.59 177.52 122.89 ;
    END
  END multdiv_ready_id_o
  PIN multdiv_signed_mode_ex_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 414.31 177.52 414.61 ;
    END
  END multdiv_signed_mode_ex_o[0]
  PIN multdiv_signed_mode_ex_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 373.51 177.52 373.81 ;
    END
  END multdiv_signed_mode_ex_o[1]
  PIN nmi_mode_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 497.95 177.52 498.25 ;
    END
  END nmi_mode_o
  PIN nt_branch_mispredict_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 79.75 0.8 80.05 ;
    END
  END nt_branch_mispredict_o
  PIN outstanding_load_wb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  174.96 0 175.1 0.485 ;
    END
  END outstanding_load_wb_i
  PIN outstanding_store_wb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  117.92 0 118.06 0.485 ;
    END
  END outstanding_store_wb_i
  PIN pc_id_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 365.35 177.52 365.65 ;
    END
  END pc_id_i[0]
  PIN pc_id_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 442.87 177.52 443.17 ;
    END
  END pc_id_i[10]
  PIN pc_id_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 432.67 177.52 432.97 ;
    END
  END pc_id_i[11]
  PIN pc_id_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 2.23 0.8 2.53 ;
    END
  END pc_id_i[12]
  PIN pc_id_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 257.23 0.8 257.53 ;
    END
  END pc_id_i[13]
  PIN pc_id_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 285.79 0.8 286.09 ;
    END
  END pc_id_i[14]
  PIN pc_id_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 291.91 0.8 292.21 ;
    END
  END pc_id_i[15]
  PIN pc_id_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 259.27 0.8 259.57 ;
    END
  END pc_id_i[16]
  PIN pc_id_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 287.83 0.8 288.13 ;
    END
  END pc_id_i[17]
  PIN pc_id_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 279.67 0.8 279.97 ;
    END
  END pc_id_i[18]
  PIN pc_id_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 198.07 0.8 198.37 ;
    END
  END pc_id_i[19]
  PIN pc_id_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 18.55 0.8 18.85 ;
    END
  END pc_id_i[1]
  PIN pc_id_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 283.75 0.8 284.05 ;
    END
  END pc_id_i[20]
  PIN pc_id_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 273.55 0.8 273.85 ;
    END
  END pc_id_i[21]
  PIN pc_id_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 240.91 0.8 241.21 ;
    END
  END pc_id_i[22]
  PIN pc_id_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 6.31 0.8 6.61 ;
    END
  END pc_id_i[23]
  PIN pc_id_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 242.95 0.8 243.25 ;
    END
  END pc_id_i[24]
  PIN pc_id_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 224.59 177.52 224.89 ;
    END
  END pc_id_i[25]
  PIN pc_id_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 214.39 177.52 214.69 ;
    END
  END pc_id_i[26]
  PIN pc_id_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 210.31 177.52 210.61 ;
    END
  END pc_id_i[27]
  PIN pc_id_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 175.63 177.52 175.93 ;
    END
  END pc_id_i[28]
  PIN pc_id_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 63.43 177.52 63.73 ;
    END
  END pc_id_i[29]
  PIN pc_id_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 128.71 177.52 129.01 ;
    END
  END pc_id_i[2]
  PIN pc_id_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 91.99 177.52 92.29 ;
    END
  END pc_id_i[30]
  PIN pc_id_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 43.03 177.52 43.33 ;
    END
  END pc_id_i[31]
  PIN pc_id_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 16.51 177.52 16.81 ;
    END
  END pc_id_i[3]
  PIN pc_id_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 2.23 177.52 2.53 ;
    END
  END pc_id_i[4]
  PIN pc_id_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 34.87 177.52 35.17 ;
    END
  END pc_id_i[5]
  PIN pc_id_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 346.99 177.52 347.29 ;
    END
  END pc_id_i[6]
  PIN pc_id_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 389.83 177.52 390.13 ;
    END
  END pc_id_i[7]
  PIN pc_id_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 422.47 177.52 422.77 ;
    END
  END pc_id_i[8]
  PIN pc_id_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 418.39 177.52 418.69 ;
    END
  END pc_id_i[9]
  PIN pc_mux_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 457.15 177.52 457.45 ;
    END
  END pc_mux_o[0]
  PIN pc_mux_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 526.51 177.52 526.81 ;
    END
  END pc_mux_o[1]
  PIN pc_mux_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 438.79 177.52 439.09 ;
    END
  END pc_mux_o[2]
  PIN pc_set_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 322.51 177.52 322.81 ;
    END
  END pc_set_o
  PIN pc_set_spec_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 324.55 177.52 324.85 ;
    END
  END pc_set_spec_o
  PIN perf_branch_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 208.27 177.52 208.57 ;
    END
  END perf_branch_o
  PIN perf_div_wait_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 120.55 177.52 120.85 ;
    END
  END perf_div_wait_o
  PIN perf_dside_wait_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 171.55 177.52 171.85 ;
    END
  END perf_dside_wait_o
  PIN perf_jump_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 179.71 177.52 180.01 ;
    END
  END perf_jump_o
  PIN perf_mul_wait_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 45.07 177.52 45.37 ;
    END
  END perf_mul_wait_o
  PIN perf_tbranch_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 489.79 177.52 490.09 ;
    END
  END perf_tbranch_o
  PIN priv_mode_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 477.55 177.52 477.85 ;
    END
  END priv_mode_i[0]
  PIN priv_mode_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 514.27 177.52 514.57 ;
    END
  END priv_mode_i[1]
  PIN ready_wb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 20.59 177.52 20.89 ;
    END
  END ready_wb_i
  PIN result_ex_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 338.83 177.52 339.13 ;
    END
  END result_ex_i[0]
  PIN result_ex_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 385.75 177.52 386.05 ;
    END
  END result_ex_i[10]
  PIN result_ex_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 430.63 177.52 430.93 ;
    END
  END result_ex_i[11]
  PIN result_ex_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 428.59 177.52 428.89 ;
    END
  END result_ex_i[12]
  PIN result_ex_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 440.83 177.52 441.13 ;
    END
  END result_ex_i[13]
  PIN result_ex_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 444.91 177.52 445.21 ;
    END
  END result_ex_i[14]
  PIN result_ex_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 434.71 177.52 435.01 ;
    END
  END result_ex_i[15]
  PIN result_ex_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 538.75 177.52 539.05 ;
    END
  END result_ex_i[16]
  PIN result_ex_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 412.27 177.52 412.57 ;
    END
  END result_ex_i[17]
  PIN result_ex_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 448.99 177.52 449.29 ;
    END
  END result_ex_i[18]
  PIN result_ex_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 495.91 177.52 496.21 ;
    END
  END result_ex_i[19]
  PIN result_ex_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 648.91 177.52 649.21 ;
    END
  END result_ex_i[1]
  PIN result_ex_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 491.83 177.52 492.13 ;
    END
  END result_ex_i[20]
  PIN result_ex_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 446.95 177.52 447.25 ;
    END
  END result_ex_i[21]
  PIN result_ex_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 485.71 177.52 486.01 ;
    END
  END result_ex_i[22]
  PIN result_ex_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 420.43 177.52 420.73 ;
    END
  END result_ex_i[23]
  PIN result_ex_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 518.35 177.52 518.65 ;
    END
  END result_ex_i[24]
  PIN result_ex_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 614.23 177.52 614.53 ;
    END
  END result_ex_i[25]
  PIN result_ex_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 453.07 177.52 453.37 ;
    END
  END result_ex_i[26]
  PIN result_ex_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 697.87 177.52 698.17 ;
    END
  END result_ex_i[27]
  PIN result_ex_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  176.72 410.23 177.52 410.53 ;
    END
  END result_ex_i[28]
  PIN result_ex_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  141.84 0 141.98 0.485 ;
    END
  END result_ex_i[29]
  PIN result_ex_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  130.8 0 130.94 0.485 ;
    END
  END result_ex_i[2]
  PIN result_ex_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  128.96 0 129.1 0.485 ;
    END
  END result_ex_i[30]
  PIN result_ex_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  140 0 140.14 0.485 ;
    END
  END result_ex_i[31]
  PIN result_ex_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  132.64 0 132.78 0.485 ;
    END
  END result_ex_i[3]
  PIN result_ex_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  138.16 0 138.3 0.485 ;
    END
  END result_ex_i[4]
  PIN result_ex_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  136.32 0 136.46 0.485 ;
    END
  END result_ex_i[5]
  PIN result_ex_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  134.48 0 134.62 0.485 ;
    END
  END result_ex_i[6]
  PIN result_ex_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  127.12 0 127.26 0.485 ;
    END
  END result_ex_i[7]
  PIN result_ex_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  119.76 0 119.9 0.485 ;
    END
  END result_ex_i[8]
  PIN result_ex_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  121.6 0 121.74 0.485 ;
    END
  END result_ex_i[9]
  PIN rf_raddr_a_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  2 703.585 2.14 704.07 ;
    END
  END rf_raddr_a_o[0]
  PIN rf_raddr_a_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  9.36 703.585 9.5 704.07 ;
    END
  END rf_raddr_a_o[1]
  PIN rf_raddr_a_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  27.76 703.585 27.9 704.07 ;
    END
  END rf_raddr_a_o[2]
  PIN rf_raddr_a_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  31.44 703.585 31.58 704.07 ;
    END
  END rf_raddr_a_o[3]
  PIN rf_raddr_a_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  40.64 703.585 40.78 704.07 ;
    END
  END rf_raddr_a_o[4]
  PIN rf_raddr_b_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  108.72 703.585 108.86 704.07 ;
    END
  END rf_raddr_b_o[0]
  PIN rf_raddr_b_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  92.16 703.585 92.3 704.07 ;
    END
  END rf_raddr_b_o[1]
  PIN rf_raddr_b_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  84.8 703.585 84.94 704.07 ;
    END
  END rf_raddr_b_o[2]
  PIN rf_raddr_b_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  88.48 703.585 88.62 704.07 ;
    END
  END rf_raddr_b_o[3]
  PIN rf_raddr_b_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  22.24 703.585 22.38 704.07 ;
    END
  END rf_raddr_b_o[4]
  PIN rf_rd_a_wb_match_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  25.92 0 26.06 0.485 ;
    END
  END rf_rd_a_wb_match_o
  PIN rf_rd_b_wb_match_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  20.4 0 20.54 0.485 ;
    END
  END rf_rd_b_wb_match_o
  PIN rf_rdata_a_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  60.88 0 61.02 0.485 ;
    END
  END rf_rdata_a_i[0]
  PIN rf_rdata_a_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  3.84 703.585 3.98 704.07 ;
    END
  END rf_rdata_a_i[10]
  PIN rf_rdata_a_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  24.08 703.585 24.22 704.07 ;
    END
  END rf_rdata_a_i[11]
  PIN rf_rdata_a_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  13.04 703.585 13.18 704.07 ;
    END
  END rf_rdata_a_i[12]
  PIN rf_rdata_a_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  20.4 703.585 20.54 704.07 ;
    END
  END rf_rdata_a_i[13]
  PIN rf_rdata_a_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  14.88 703.585 15.02 704.07 ;
    END
  END rf_rdata_a_i[14]
  PIN rf_rdata_a_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  18.56 703.585 18.7 704.07 ;
    END
  END rf_rdata_a_i[15]
  PIN rf_rdata_a_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  16.72 703.585 16.86 704.07 ;
    END
  END rf_rdata_a_i[16]
  PIN rf_rdata_a_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  36.96 703.585 37.1 704.07 ;
    END
  END rf_rdata_a_i[17]
  PIN rf_rdata_a_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  18.56 0 18.7 0.485 ;
    END
  END rf_rdata_a_i[18]
  PIN rf_rdata_a_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  42.48 0 42.62 0.485 ;
    END
  END rf_rdata_a_i[19]
  PIN rf_rdata_a_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  53.52 0 53.66 0.485 ;
    END
  END rf_rdata_a_i[1]
  PIN rf_rdata_a_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  22.24 0 22.38 0.485 ;
    END
  END rf_rdata_a_i[20]
  PIN rf_rdata_a_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  27.76 0 27.9 0.485 ;
    END
  END rf_rdata_a_i[21]
  PIN rf_rdata_a_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  44.32 0 44.46 0.485 ;
    END
  END rf_rdata_a_i[22]
  PIN rf_rdata_a_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  40.64 0 40.78 0.485 ;
    END
  END rf_rdata_a_i[23]
  PIN rf_rdata_a_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  24.08 0 24.22 0.485 ;
    END
  END rf_rdata_a_i[24]
  PIN rf_rdata_a_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  29.6 0 29.74 0.485 ;
    END
  END rf_rdata_a_i[25]
  PIN rf_rdata_a_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  35.12 0 35.26 0.485 ;
    END
  END rf_rdata_a_i[26]
  PIN rf_rdata_a_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  38.8 0 38.94 0.485 ;
    END
  END rf_rdata_a_i[27]
  PIN rf_rdata_a_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  46.16 0 46.3 0.485 ;
    END
  END rf_rdata_a_i[28]
  PIN rf_rdata_a_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  49.84 0 49.98 0.485 ;
    END
  END rf_rdata_a_i[29]
  PIN rf_rdata_a_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  59.04 0 59.18 0.485 ;
    END
  END rf_rdata_a_i[2]
  PIN rf_rdata_a_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  55.36 0 55.5 0.485 ;
    END
  END rf_rdata_a_i[30]
  PIN rf_rdata_a_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  64.56 0 64.7 0.485 ;
    END
  END rf_rdata_a_i[31]
  PIN rf_rdata_a_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  57.2 0 57.34 0.485 ;
    END
  END rf_rdata_a_i[3]
  PIN rf_rdata_a_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  51.68 0 51.82 0.485 ;
    END
  END rf_rdata_a_i[4]
  PIN rf_rdata_a_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  66.4 0 66.54 0.485 ;
    END
  END rf_rdata_a_i[5]
  PIN rf_rdata_a_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  62.72 0 62.86 0.485 ;
    END
  END rf_rdata_a_i[6]
  PIN rf_rdata_a_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  57.2 703.585 57.34 704.07 ;
    END
  END rf_rdata_a_i[7]
  PIN rf_rdata_a_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  51.68 703.585 51.82 704.07 ;
    END
  END rf_rdata_a_i[8]
  PIN rf_rdata_a_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  103.2 703.585 103.34 704.07 ;
    END
  END rf_rdata_a_i[9]
  PIN rf_rdata_b_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  95.84 703.585 95.98 704.07 ;
    END
  END rf_rdata_b_i[0]
  PIN rf_rdata_b_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  81.12 703.585 81.26 704.07 ;
    END
  END rf_rdata_b_i[10]
  PIN rf_rdata_b_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  105.04 703.585 105.18 704.07 ;
    END
  END rf_rdata_b_i[11]
  PIN rf_rdata_b_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  44.32 703.585 44.46 704.07 ;
    END
  END rf_rdata_b_i[12]
  PIN rf_rdata_b_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  7.52 703.585 7.66 704.07 ;
    END
  END rf_rdata_b_i[13]
  PIN rf_rdata_b_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  48 703.585 48.14 704.07 ;
    END
  END rf_rdata_b_i[14]
  PIN rf_rdata_b_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  29.6 703.585 29.74 704.07 ;
    END
  END rf_rdata_b_i[15]
  PIN rf_rdata_b_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  5.68 703.585 5.82 704.07 ;
    END
  END rf_rdata_b_i[16]
  PIN rf_rdata_b_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  33.28 703.585 33.42 704.07 ;
    END
  END rf_rdata_b_i[17]
  PIN rf_rdata_b_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  25.92 703.585 26.06 704.07 ;
    END
  END rf_rdata_b_i[18]
  PIN rf_rdata_b_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  46.16 703.585 46.3 704.07 ;
    END
  END rf_rdata_b_i[19]
  PIN rf_rdata_b_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  53.52 703.585 53.66 704.07 ;
    END
  END rf_rdata_b_i[1]
  PIN rf_rdata_b_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  49.84 703.585 49.98 704.07 ;
    END
  END rf_rdata_b_i[20]
  PIN rf_rdata_b_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  35.12 703.585 35.26 704.07 ;
    END
  END rf_rdata_b_i[21]
  PIN rf_rdata_b_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  59.04 703.585 59.18 704.07 ;
    END
  END rf_rdata_b_i[22]
  PIN rf_rdata_b_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  11.2 703.585 11.34 704.07 ;
    END
  END rf_rdata_b_i[23]
  PIN rf_rdata_b_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  42.48 703.585 42.62 704.07 ;
    END
  END rf_rdata_b_i[24]
  PIN rf_rdata_b_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  66.4 703.585 66.54 704.07 ;
    END
  END rf_rdata_b_i[25]
  PIN rf_rdata_b_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  99.52 703.585 99.66 704.07 ;
    END
  END rf_rdata_b_i[26]
  PIN rf_rdata_b_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  71.92 703.585 72.06 704.07 ;
    END
  END rf_rdata_b_i[27]
  PIN rf_rdata_b_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  97.68 703.585 97.82 704.07 ;
    END
  END rf_rdata_b_i[28]
  PIN rf_rdata_b_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  75.6 703.585 75.74 704.07 ;
    END
  END rf_rdata_b_i[29]
  PIN rf_rdata_b_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  106.88 703.585 107.02 704.07 ;
    END
  END rf_rdata_b_i[2]
  PIN rf_rdata_b_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  70.08 703.585 70.22 704.07 ;
    END
  END rf_rdata_b_i[30]
  PIN rf_rdata_b_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  64.56 703.585 64.7 704.07 ;
    END
  END rf_rdata_b_i[31]
  PIN rf_rdata_b_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  62.72 703.585 62.86 704.07 ;
    END
  END rf_rdata_b_i[3]
  PIN rf_rdata_b_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  55.36 703.585 55.5 704.07 ;
    END
  END rf_rdata_b_i[4]
  PIN rf_rdata_b_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  77.44 703.585 77.58 704.07 ;
    END
  END rf_rdata_b_i[5]
  PIN rf_rdata_b_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  90.32 703.585 90.46 704.07 ;
    END
  END rf_rdata_b_i[6]
  PIN rf_rdata_b_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  94 703.585 94.14 704.07 ;
    END
  END rf_rdata_b_i[7]
  PIN rf_rdata_b_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  82.96 703.585 83.1 704.07 ;
    END
  END rf_rdata_b_i[8]
  PIN rf_rdata_b_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  86.64 703.585 86.78 704.07 ;
    END
  END rf_rdata_b_i[9]
  PIN rf_ren_a_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  81.12 0 81.26 0.485 ;
    END
  END rf_ren_a_o
  PIN rf_ren_b_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  82.96 0 83.1 0.485 ;
    END
  END rf_ren_b_o
  PIN rf_waddr_id_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  79.28 703.585 79.42 704.07 ;
    END
  END rf_waddr_id_o[0]
  PIN rf_waddr_id_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  60.88 703.585 61.02 704.07 ;
    END
  END rf_waddr_id_o[1]
  PIN rf_waddr_id_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  73.76 703.585 73.9 704.07 ;
    END
  END rf_waddr_id_o[2]
  PIN rf_waddr_id_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  68.24 703.585 68.38 704.07 ;
    END
  END rf_waddr_id_o[3]
  PIN rf_waddr_id_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  38.8 703.585 38.94 704.07 ;
    END
  END rf_waddr_id_o[4]
  PIN rf_waddr_wb_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  169.44 0 169.58 0.485 ;
    END
  END rf_waddr_wb_i[0]
  PIN rf_waddr_wb_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  105.04 0 105.18 0.485 ;
    END
  END rf_waddr_wb_i[1]
  PIN rf_waddr_wb_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  101.36 0 101.5 0.485 ;
    END
  END rf_waddr_wb_i[2]
  PIN rf_waddr_wb_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  33.28 0 33.42 0.485 ;
    END
  END rf_waddr_wb_i[3]
  PIN rf_waddr_wb_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  11.2 0 11.34 0.485 ;
    END
  END rf_waddr_wb_i[4]
  PIN rf_wdata_fwd_wb_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  147.36 0 147.5 0.485 ;
    END
  END rf_wdata_fwd_wb_i[0]
  PIN rf_wdata_fwd_wb_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  86.64 0 86.78 0.485 ;
    END
  END rf_wdata_fwd_wb_i[10]
  PIN rf_wdata_fwd_wb_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  167.6 0 167.74 0.485 ;
    END
  END rf_wdata_fwd_wb_i[11]
  PIN rf_wdata_fwd_wb_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  163.92 0 164.06 0.485 ;
    END
  END rf_wdata_fwd_wb_i[12]
  PIN rf_wdata_fwd_wb_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  112.4 0 112.54 0.485 ;
    END
  END rf_wdata_fwd_wb_i[13]
  PIN rf_wdata_fwd_wb_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  88.48 0 88.62 0.485 ;
    END
  END rf_wdata_fwd_wb_i[14]
  PIN rf_wdata_fwd_wb_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  103.2 0 103.34 0.485 ;
    END
  END rf_wdata_fwd_wb_i[15]
  PIN rf_wdata_fwd_wb_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  156.56 0 156.7 0.485 ;
    END
  END rf_wdata_fwd_wb_i[16]
  PIN rf_wdata_fwd_wb_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  68.24 0 68.38 0.485 ;
    END
  END rf_wdata_fwd_wb_i[17]
  PIN rf_wdata_fwd_wb_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  36.96 0 37.1 0.485 ;
    END
  END rf_wdata_fwd_wb_i[18]
  PIN rf_wdata_fwd_wb_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  70.08 0 70.22 0.485 ;
    END
  END rf_wdata_fwd_wb_i[19]
  PIN rf_wdata_fwd_wb_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  73.76 0 73.9 0.485 ;
    END
  END rf_wdata_fwd_wb_i[1]
  PIN rf_wdata_fwd_wb_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  84.8 0 84.94 0.485 ;
    END
  END rf_wdata_fwd_wb_i[20]
  PIN rf_wdata_fwd_wb_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  149.2 0 149.34 0.485 ;
    END
  END rf_wdata_fwd_wb_i[21]
  PIN rf_wdata_fwd_wb_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  77.44 0 77.58 0.485 ;
    END
  END rf_wdata_fwd_wb_i[22]
  PIN rf_wdata_fwd_wb_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  16.72 0 16.86 0.485 ;
    END
  END rf_wdata_fwd_wb_i[23]
  PIN rf_wdata_fwd_wb_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  92.16 0 92.3 0.485 ;
    END
  END rf_wdata_fwd_wb_i[24]
  PIN rf_wdata_fwd_wb_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  79.28 0 79.42 0.485 ;
    END
  END rf_wdata_fwd_wb_i[25]
  PIN rf_wdata_fwd_wb_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  114.24 0 114.38 0.485 ;
    END
  END rf_wdata_fwd_wb_i[26]
  PIN rf_wdata_fwd_wb_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  31.44 0 31.58 0.485 ;
    END
  END rf_wdata_fwd_wb_i[27]
  PIN rf_wdata_fwd_wb_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  90.32 0 90.46 0.485 ;
    END
  END rf_wdata_fwd_wb_i[28]
  PIN rf_wdata_fwd_wb_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  116.08 0 116.22 0.485 ;
    END
  END rf_wdata_fwd_wb_i[29]
  PIN rf_wdata_fwd_wb_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  7.52 0 7.66 0.485 ;
    END
  END rf_wdata_fwd_wb_i[2]
  PIN rf_wdata_fwd_wb_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  95.84 0 95.98 0.485 ;
    END
  END rf_wdata_fwd_wb_i[30]
  PIN rf_wdata_fwd_wb_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  97.68 0 97.82 0.485 ;
    END
  END rf_wdata_fwd_wb_i[31]
  PIN rf_wdata_fwd_wb_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  171.28 0 171.42 0.485 ;
    END
  END rf_wdata_fwd_wb_i[3]
  PIN rf_wdata_fwd_wb_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  99.52 0 99.66 0.485 ;
    END
  END rf_wdata_fwd_wb_i[4]
  PIN rf_wdata_fwd_wb_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  151.04 0 151.18 0.485 ;
    END
  END rf_wdata_fwd_wb_i[5]
  PIN rf_wdata_fwd_wb_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  14.88 0 15.02 0.485 ;
    END
  END rf_wdata_fwd_wb_i[6]
  PIN rf_wdata_fwd_wb_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  165.76 0 165.9 0.485 ;
    END
  END rf_wdata_fwd_wb_i[7]
  PIN rf_wdata_fwd_wb_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  106.88 0 107.02 0.485 ;
    END
  END rf_wdata_fwd_wb_i[8]
  PIN rf_wdata_fwd_wb_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  110.56 0 110.7 0.485 ;
    END
  END rf_wdata_fwd_wb_i[9]
  PIN rf_wdata_id_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  125.28 0 125.42 0.485 ;
    END
  END rf_wdata_id_o[0]
  PIN rf_wdata_id_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  123.44 0 123.58 0.485 ;
    END
  END rf_wdata_id_o[10]
  PIN rf_wdata_id_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  121.6 703.585 121.74 704.07 ;
    END
  END rf_wdata_id_o[11]
  PIN rf_wdata_id_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  114.24 703.585 114.38 704.07 ;
    END
  END rf_wdata_id_o[12]
  PIN rf_wdata_id_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  123.44 703.585 123.58 704.07 ;
    END
  END rf_wdata_id_o[13]
  PIN rf_wdata_id_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  125.28 703.585 125.42 704.07 ;
    END
  END rf_wdata_id_o[14]
  PIN rf_wdata_id_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  112.4 703.585 112.54 704.07 ;
    END
  END rf_wdata_id_o[15]
  PIN rf_wdata_id_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  117.92 703.585 118.06 704.07 ;
    END
  END rf_wdata_id_o[16]
  PIN rf_wdata_id_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  116.08 703.585 116.22 704.07 ;
    END
  END rf_wdata_id_o[17]
  PIN rf_wdata_id_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  165.76 703.585 165.9 704.07 ;
    END
  END rf_wdata_id_o[18]
  PIN rf_wdata_id_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  160.24 703.585 160.38 704.07 ;
    END
  END rf_wdata_id_o[19]
  PIN rf_wdata_id_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  143.68 703.585 143.82 704.07 ;
    END
  END rf_wdata_id_o[1]
  PIN rf_wdata_id_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  152.88 703.585 153.02 704.07 ;
    END
  END rf_wdata_id_o[20]
  PIN rf_wdata_id_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  151.04 703.585 151.18 704.07 ;
    END
  END rf_wdata_id_o[21]
  PIN rf_wdata_id_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  138.16 703.585 138.3 704.07 ;
    END
  END rf_wdata_id_o[22]
  PIN rf_wdata_id_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  145.52 703.585 145.66 704.07 ;
    END
  END rf_wdata_id_o[23]
  PIN rf_wdata_id_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  134.48 703.585 134.62 704.07 ;
    END
  END rf_wdata_id_o[24]
  PIN rf_wdata_id_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  147.36 703.585 147.5 704.07 ;
    END
  END rf_wdata_id_o[25]
  PIN rf_wdata_id_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  149.2 703.585 149.34 704.07 ;
    END
  END rf_wdata_id_o[26]
  PIN rf_wdata_id_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  140 703.585 140.14 704.07 ;
    END
  END rf_wdata_id_o[27]
  PIN rf_wdata_id_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  163.92 703.585 164.06 704.07 ;
    END
  END rf_wdata_id_o[28]
  PIN rf_wdata_id_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  158.4 703.585 158.54 704.07 ;
    END
  END rf_wdata_id_o[29]
  PIN rf_wdata_id_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  130.8 703.585 130.94 704.07 ;
    END
  END rf_wdata_id_o[2]
  PIN rf_wdata_id_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  162.08 703.585 162.22 704.07 ;
    END
  END rf_wdata_id_o[30]
  PIN rf_wdata_id_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  154.72 703.585 154.86 704.07 ;
    END
  END rf_wdata_id_o[31]
  PIN rf_wdata_id_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  132.64 703.585 132.78 704.07 ;
    END
  END rf_wdata_id_o[3]
  PIN rf_wdata_id_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  156.56 703.585 156.7 704.07 ;
    END
  END rf_wdata_id_o[4]
  PIN rf_wdata_id_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  136.32 703.585 136.46 704.07 ;
    END
  END rf_wdata_id_o[5]
  PIN rf_wdata_id_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  141.84 703.585 141.98 704.07 ;
    END
  END rf_wdata_id_o[6]
  PIN rf_wdata_id_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  128.96 703.585 129.1 704.07 ;
    END
  END rf_wdata_id_o[7]
  PIN rf_wdata_id_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  119.76 703.585 119.9 704.07 ;
    END
  END rf_wdata_id_o[8]
  PIN rf_wdata_id_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  110.56 703.585 110.7 704.07 ;
    END
  END rf_wdata_id_o[9]
  PIN rf_we_id_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  101.36 703.585 101.5 704.07 ;
    END
  END rf_we_id_o
  PIN rf_write_wb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  174.96 703.585 175.1 704.07 ;
    END
  END rf_write_wb_i
  PIN rst_ni
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  171.28 703.585 171.42 704.07 ;
    END
  END rst_ni
  PIN trigger_match_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  127.12 703.585 127.26 704.07 ;
    END
  END trigger_match_i
  OBS
    LAYER nwell ;
     RECT  0 0 177.52 704.07 ;
    LAYER pwell ;
     RECT  0 0 177.52 704.07 ;
    LAYER li1 ;
     RECT  0 0 177.52 704.07 ;
    LAYER met1 ;
     RECT  0 0 177.52 704.07 ;
    LAYER met2 ;
     RECT  0 0 177.52 704.07 ;
    LAYER met3 ;
     RECT  0 0 177.52 704.07 ;
    LAYER met4 ;
     RECT  0 0 177.52 704.07 ;
    LAYER met5 ;
     RECT  0 0 177.52 704.07 ;
  END
END ibex_id_stage
END LIBRARY
